`ifdef ST_WIDTH_INF_4
reg [63:0] gol_yjp0  ;
reg [63:0] gol_yjp1  ;
reg [63:0] dut_yjp0  ;
reg [63:0] dut_yjp1  ;
`endif //ST_WIDTH_INF_4
`ifdef ST_WIDTH_INF_4
real gol_re_yjp0  ;
real gol_re_yjp1  ;
real gol_im_yjp0  ;
real gol_im_yjp1  ;
real dut_re_yjp0  ;
real dut_re_yjp1  ;
real dut_im_yjp0  ;
real dut_im_yjp1  ;
`endif //ST_WIDTH_INF_4
`ifdef ST_WIDTH_INF_4
real err_re_per0   ;    
real err_re_per1   ;    
real err_im_per0   ;    
real err_im_per1   ;    
`endif //ST_WIDTH_INF_4

`ifdef ST_WIDTH_INF_8
reg [63:0] gol_yjp0  ;
reg [63:0] gol_yjp1  ;
reg [63:0] dut_yjp0  ;
reg [63:0] dut_yjp1  ;
reg [63:0] gol_yjp2  ;
reg [63:0] gol_yjp3  ;
reg [63:0] dut_yjp2  ;
reg [63:0] dut_yjp3  ;

`endif //ST_WIDTH_INF_8
`ifdef ST_WIDTH_INF_8
real gol_re_yjp0  ;
real gol_re_yjp1  ;
real gol_im_yjp0  ;
real gol_im_yjp1  ;
real dut_re_yjp0  ;
real dut_re_yjp1  ;
real dut_im_yjp0  ;
real dut_im_yjp1  ;
//
real gol_re_yjp2  ;
real gol_re_yjp3  ;
real gol_im_yjp2  ;
real gol_im_yjp3  ;
real dut_re_yjp2  ;
real dut_re_yjp3  ;
real dut_im_yjp2  ;
real dut_im_yjp3  ;

`endif //ST_WIDTH_INF_8
`ifdef ST_WIDTH_INF_8
real err_re_per0   ;    
real err_re_per1   ;    
real err_im_per0   ;    
real err_im_per1   ;
real err_re_per2   ;    
real err_re_per3   ;    
real err_im_per2   ;    
real err_im_per3   ; 
`endif //ST_WIDTH_INF_4
