`ifdef ST_WIDTH_INF_4
$fwrite(tri_report, "===============================%d Column Results    ======================================\n",col_index);
if(col_index>=0  ) begin if(err_re_per0  <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item0 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per0  , gol_re_yjp0  , dut_re_yjp0  ); end else begin $fwrite(tri_report, "Item0 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per0  , gol_re_yjp0  , dut_re_yjp0  ); end end
if(col_index>=0  ) begin if(err_im_per0  <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item0 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per0  , gol_im_yjp0  , dut_im_yjp0  ); end else begin $fwrite(tri_report, "Item0 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per0  , gol_im_yjp0  , dut_im_yjp0  ); end end

if(col_index>=1  ) begin if(err_re_per1  <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item1 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per1  , gol_re_yjp1  , dut_re_yjp1  ); end else begin $fwrite(tri_report, "Item1 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per1  , gol_re_yjp1  , dut_re_yjp1  ); end end
if(col_index>=1  ) begin if(err_im_per1  <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item1 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per1  , gol_im_yjp1  , dut_im_yjp1  ); end else begin $fwrite(tri_report, "Item1 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per1  , gol_im_yjp1  , dut_im_yjp1  ); end end
`endif // ST_WIDTH_INF_4
