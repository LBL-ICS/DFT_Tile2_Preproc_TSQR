`ifdef ST_WIDTH_INF_4
reg [63:0] gol_yjp0  ;
reg [63:0] gol_yjp1  ;
reg [63:0] dut_yjp0  ;
reg [63:0] dut_yjp1  ;
`endif //ST_WIDTH_INF_4
`ifdef ST_WIDTH_INF_4
real gol_re_yjp0  ;
real gol_re_yjp1  ;
real gol_im_yjp0  ;
real gol_im_yjp1  ;
real dut_re_yjp0  ;
real dut_re_yjp1  ;
real dut_im_yjp0  ;
real dut_im_yjp1  ;
`endif //ST_WIDTH_INF_4
`ifdef ST_WIDTH_INF_4
real err_re_per0   ;    
real err_re_per1   ;    
real err_im_per0   ;    
real err_im_per1   ;    
`endif //ST_WIDTH_INF_4
