`ifdef ST_WIDTH_INF_4
$fwrite(tri_report, "===============================%d Column Results    ======================================\n",col_index);
if(col_index>=0  ) begin if(err_re_per0  <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item0 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per0  , gol_re_yjp0  , dut_re_yjp0  ); end else begin $fwrite(tri_report, "Item0 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per0  , gol_re_yjp0  , dut_re_yjp0  ); end end
if(col_index>=0  ) begin if(err_im_per0  <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item0 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per0  , gol_im_yjp0  , dut_im_yjp0  ); end else begin $fwrite(tri_report, "Item0 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per0  , gol_im_yjp0  , dut_im_yjp0  ); end end

if(col_index>=1  ) begin if(err_re_per1  <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item1 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per1  , gol_re_yjp1  , dut_re_yjp1  ); end else begin $fwrite(tri_report, "Item1 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per1  , gol_re_yjp1  , dut_re_yjp1  ); end end
if(col_index>=1  ) begin if(err_im_per1  <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item1 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per1  , gol_im_yjp1  , dut_im_yjp1  ); end else begin $fwrite(tri_report, "Item1 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per1  , gol_im_yjp1  , dut_im_yjp1  ); end end
`endif // ST_WIDTH_INF_4


`ifdef ST_WIDTH_INF_8
$fwrite(tri_report, "===============================%d Column Results    ======================================\n",col_index);
if(col_index>=0  ) begin if(err_re_per0  <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item0 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per0  , gol_re_yjp0  , dut_re_yjp0  ); end else begin $fwrite(tri_report, "Item0 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per0  , gol_re_yjp0  , dut_re_yjp0  ); end end
if(col_index>=0  ) begin if(err_im_per0  <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item0 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per0  , gol_im_yjp0  , dut_im_yjp0  ); end else begin $fwrite(tri_report, "Item0 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per0  , gol_im_yjp0  , dut_im_yjp0  ); end end

if(col_index>=1  ) begin if(err_re_per1  <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item1 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per1  , gol_re_yjp1  , dut_re_yjp1  ); end else begin $fwrite(tri_report, "Item1 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per1  , gol_re_yjp1  , dut_re_yjp1  ); end end
if(col_index>=1  ) begin if(err_im_per1  <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item1 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per1  , gol_im_yjp1  , dut_im_yjp1  ); end else begin $fwrite(tri_report, "Item1 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per1  , gol_im_yjp1  , dut_im_yjp1  ); end end
//
if(col_index>=2  ) begin if(err_re_per2  <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item2 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per2  , gol_re_yjp2  , dut_re_yjp2  ); end else begin $fwrite(tri_report, "Item0 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per2  , gol_re_yjp2  , dut_re_yjp2  ); end end
if(col_index>=2  ) begin if(err_im_per2  <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item2 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per2  , gol_im_yjp2  , dut_im_yjp2  ); end else begin $fwrite(tri_report, "Item0 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per2  , gol_im_yjp2  , dut_im_yjp2  ); end end

if(col_index>=3  ) begin if(err_re_per3  <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item3 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per3  , gol_re_yjp3  , dut_re_yjp3  ); end else begin $fwrite(tri_report, "Item3 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per3  , gol_re_yjp3  , dut_re_yjp3  ); end end
if(col_index>=3  ) begin if(err_im_per3  <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item3 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per3  , gol_im_yjp3  , dut_im_yjp3  ); end else begin $fwrite(tri_report, "Item3 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per3  , gol_im_yjp3  , dut_im_yjp3  ); end end

`endif // ST_WIDTH_INF_4


`ifdef ST_WIDTH_INF_16
if(col_index>=0) begin if(err_re_per0 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item0 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per0, gol_re_yjp0, dut_re_yjp0); end else begin $fwrite(tri_report, "Item0 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per0, gol_re_yjp0, dut_re_yjp0); end end
if(col_index>=0) begin if(err_im_per0 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item0 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per0, gol_im_yjp0, dut_im_yjp0); end else begin $fwrite(tri_report, "Item0 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per0, gol_im_yjp0, dut_im_yjp0); end end

if(col_index>=1) begin if(err_re_per1 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item1 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per1, gol_re_yjp1, dut_re_yjp1); end else begin $fwrite(tri_report, "Item1 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per1, gol_re_yjp1, dut_re_yjp1); end end
if(col_index>=1) begin if(err_im_per1 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item1 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per1, gol_im_yjp1, dut_im_yjp1); end else begin $fwrite(tri_report, "Item1 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per1, gol_im_yjp1, dut_im_yjp1); end end

if(col_index>=2) begin if(err_re_per2 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item2 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per2, gol_re_yjp2, dut_re_yjp2); end else begin $fwrite(tri_report, "Item2 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per2, gol_re_yjp2, dut_re_yjp2); end end
if(col_index>=2) begin if(err_im_per2 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item2 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per2, gol_im_yjp2, dut_im_yjp2); end else begin $fwrite(tri_report, "Item2 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per2, gol_im_yjp2, dut_im_yjp2); end end

if(col_index>=3) begin if(err_re_per3 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item3 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per3, gol_re_yjp3, dut_re_yjp3); end else begin $fwrite(tri_report, "Item3 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per3, gol_re_yjp3, dut_re_yjp3); end end
if(col_index>=3) begin if(err_im_per3 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item3 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per3, gol_im_yjp3, dut_im_yjp3); end else begin $fwrite(tri_report, "Item3 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per3, gol_im_yjp3, dut_im_yjp3); end end

if(col_index>=4) begin if(err_re_per4 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item4 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per4, gol_re_yjp4, dut_re_yjp4); end else begin $fwrite(tri_report, "Item4 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per4, gol_re_yjp4, dut_re_yjp4); end end
if(col_index>=4) begin if(err_im_per4 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item4 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per4, gol_im_yjp4, dut_im_yjp4); end else begin $fwrite(tri_report, "Item4 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per4, gol_im_yjp4, dut_im_yjp4); end end

if(col_index>=5) begin if(err_re_per5 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item5 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per5, gol_re_yjp5, dut_re_yjp5); end else begin $fwrite(tri_report, "Item5 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per5, gol_re_yjp5, dut_re_yjp5); end end
if(col_index>=5) begin if(err_im_per5 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item5 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per5, gol_im_yjp5, dut_im_yjp5); end else begin $fwrite(tri_report, "Item5 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per5, gol_im_yjp5, dut_im_yjp5); end end

if(col_index>=6) begin if(err_re_per6 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item6 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per6, gol_re_yjp6, dut_re_yjp6); end else begin $fwrite(tri_report, "Item6 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per6, gol_re_yjp6, dut_re_yjp6); end end
if(col_index>=6) begin if(err_im_per6 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item6 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per6, gol_im_yjp6, dut_im_yjp6); end else begin $fwrite(tri_report, "Item6 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per6, gol_im_yjp6, dut_im_yjp6); end end

if(col_index>=7) begin if(err_re_per7 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item7 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per7, gol_re_yjp7, dut_re_yjp7); end else begin $fwrite(tri_report, "Item7 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per7, gol_re_yjp7, dut_re_yjp7); end end
if(col_index>=7) begin if(err_im_per7 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item7 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per7, gol_im_yjp7, dut_im_yjp7); end else begin $fwrite(tri_report, "Item7 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per7, gol_im_yjp7, dut_im_yjp7); end end

`endif


`ifdef ST_WIDTH_INF_512
if(col_index>=0) begin if(err_re_per0 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item0 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per0, gol_re_yjp0, dut_re_yjp0); end else begin $fwrite(tri_report, "Item0 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per0, gol_re_yjp0, dut_re_yjp0); end end
if(col_index>=0) begin if(err_im_per0 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item0 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per0, gol_im_yjp0, dut_im_yjp0); end else begin $fwrite(tri_report, "Item0 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per0, gol_im_yjp0, dut_im_yjp0); end end

if(col_index>=1) begin if(err_re_per1 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item1 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per1, gol_re_yjp1, dut_re_yjp1); end else begin $fwrite(tri_report, "Item1 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per1, gol_re_yjp1, dut_re_yjp1); end end
if(col_index>=1) begin if(err_im_per1 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item1 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per1, gol_im_yjp1, dut_im_yjp1); end else begin $fwrite(tri_report, "Item1 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per1, gol_im_yjp1, dut_im_yjp1); end end

if(col_index>=2) begin if(err_re_per2 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item2 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per2, gol_re_yjp2, dut_re_yjp2); end else begin $fwrite(tri_report, "Item2 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per2, gol_re_yjp2, dut_re_yjp2); end end
if(col_index>=2) begin if(err_im_per2 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item2 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per2, gol_im_yjp2, dut_im_yjp2); end else begin $fwrite(tri_report, "Item2 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per2, gol_im_yjp2, dut_im_yjp2); end end

if(col_index>=3) begin if(err_re_per3 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item3 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per3, gol_re_yjp3, dut_re_yjp3); end else begin $fwrite(tri_report, "Item3 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per3, gol_re_yjp3, dut_re_yjp3); end end
if(col_index>=3) begin if(err_im_per3 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item3 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per3, gol_im_yjp3, dut_im_yjp3); end else begin $fwrite(tri_report, "Item3 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per3, gol_im_yjp3, dut_im_yjp3); end end

if(col_index>=4) begin if(err_re_per4 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item4 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per4, gol_re_yjp4, dut_re_yjp4); end else begin $fwrite(tri_report, "Item4 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per4, gol_re_yjp4, dut_re_yjp4); end end
if(col_index>=4) begin if(err_im_per4 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item4 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per4, gol_im_yjp4, dut_im_yjp4); end else begin $fwrite(tri_report, "Item4 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per4, gol_im_yjp4, dut_im_yjp4); end end

if(col_index>=5) begin if(err_re_per5 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item5 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per5, gol_re_yjp5, dut_re_yjp5); end else begin $fwrite(tri_report, "Item5 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per5, gol_re_yjp5, dut_re_yjp5); end end
if(col_index>=5) begin if(err_im_per5 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item5 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per5, gol_im_yjp5, dut_im_yjp5); end else begin $fwrite(tri_report, "Item5 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per5, gol_im_yjp5, dut_im_yjp5); end end

if(col_index>=6) begin if(err_re_per6 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item6 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per6, gol_re_yjp6, dut_re_yjp6); end else begin $fwrite(tri_report, "Item6 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per6, gol_re_yjp6, dut_re_yjp6); end end
if(col_index>=6) begin if(err_im_per6 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item6 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per6, gol_im_yjp6, dut_im_yjp6); end else begin $fwrite(tri_report, "Item6 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per6, gol_im_yjp6, dut_im_yjp6); end end

if(col_index>=7) begin if(err_re_per7 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item7 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per7, gol_re_yjp7, dut_re_yjp7); end else begin $fwrite(tri_report, "Item7 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per7, gol_re_yjp7, dut_re_yjp7); end end
if(col_index>=7) begin if(err_im_per7 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item7 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per7, gol_im_yjp7, dut_im_yjp7); end else begin $fwrite(tri_report, "Item7 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per7, gol_im_yjp7, dut_im_yjp7); end end

if(col_index>=8) begin if(err_re_per8 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item8 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per8, gol_re_yjp8, dut_re_yjp8); end else begin $fwrite(tri_report, "Item8 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per8, gol_re_yjp8, dut_re_yjp8); end end
if(col_index>=8) begin if(err_im_per8 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item8 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per8, gol_im_yjp8, dut_im_yjp8); end else begin $fwrite(tri_report, "Item8 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per8, gol_im_yjp8, dut_im_yjp8); end end

if(col_index>=9) begin if(err_re_per9 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item9 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per9, gol_re_yjp9, dut_re_yjp9); end else begin $fwrite(tri_report, "Item9 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per9, gol_re_yjp9, dut_re_yjp9); end end
if(col_index>=9) begin if(err_im_per9 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item9 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per9, gol_im_yjp9, dut_im_yjp9); end else begin $fwrite(tri_report, "Item9 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per9, gol_im_yjp9, dut_im_yjp9); end end

if(col_index>=10) begin if(err_re_per10 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item10 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per10, gol_re_yjp10, dut_re_yjp10); end else begin $fwrite(tri_report, "Item10 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per10, gol_re_yjp10, dut_re_yjp10); end end
if(col_index>=10) begin if(err_im_per10 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item10 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per10, gol_im_yjp10, dut_im_yjp10); end else begin $fwrite(tri_report, "Item10 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per10, gol_im_yjp10, dut_im_yjp10); end end

if(col_index>=11) begin if(err_re_per11 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item11 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per11, gol_re_yjp11, dut_re_yjp11); end else begin $fwrite(tri_report, "Item11 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per11, gol_re_yjp11, dut_re_yjp11); end end
if(col_index>=11) begin if(err_im_per11 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item11 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per11, gol_im_yjp11, dut_im_yjp11); end else begin $fwrite(tri_report, "Item11 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per11, gol_im_yjp11, dut_im_yjp11); end end

if(col_index>=12) begin if(err_re_per12 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item12 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per12, gol_re_yjp12, dut_re_yjp12); end else begin $fwrite(tri_report, "Item12 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per12, gol_re_yjp12, dut_re_yjp12); end end
if(col_index>=12) begin if(err_im_per12 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item12 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per12, gol_im_yjp12, dut_im_yjp12); end else begin $fwrite(tri_report, "Item12 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per12, gol_im_yjp12, dut_im_yjp12); end end

if(col_index>=13) begin if(err_re_per13 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item13 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per13, gol_re_yjp13, dut_re_yjp13); end else begin $fwrite(tri_report, "Item13 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per13, gol_re_yjp13, dut_re_yjp13); end end
if(col_index>=13) begin if(err_im_per13 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item13 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per13, gol_im_yjp13, dut_im_yjp13); end else begin $fwrite(tri_report, "Item13 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per13, gol_im_yjp13, dut_im_yjp13); end end

if(col_index>=14) begin if(err_re_per14 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item14 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per14, gol_re_yjp14, dut_re_yjp14); end else begin $fwrite(tri_report, "Item14 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per14, gol_re_yjp14, dut_re_yjp14); end end
if(col_index>=14) begin if(err_im_per14 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item14 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per14, gol_im_yjp14, dut_im_yjp14); end else begin $fwrite(tri_report, "Item14 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per14, gol_im_yjp14, dut_im_yjp14); end end

if(col_index>=15) begin if(err_re_per15 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item15 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per15, gol_re_yjp15, dut_re_yjp15); end else begin $fwrite(tri_report, "Item15 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per15, gol_re_yjp15, dut_re_yjp15); end end
if(col_index>=15) begin if(err_im_per15 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item15 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per15, gol_im_yjp15, dut_im_yjp15); end else begin $fwrite(tri_report, "Item15 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per15, gol_im_yjp15, dut_im_yjp15); end end

if(col_index>=16) begin if(err_re_per16 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item16 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per16, gol_re_yjp16, dut_re_yjp16); end else begin $fwrite(tri_report, "Item16 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per16, gol_re_yjp16, dut_re_yjp16); end end
if(col_index>=16) begin if(err_im_per16 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item16 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per16, gol_im_yjp16, dut_im_yjp16); end else begin $fwrite(tri_report, "Item16 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per16, gol_im_yjp16, dut_im_yjp16); end end

if(col_index>=17) begin if(err_re_per17 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item17 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per17, gol_re_yjp17, dut_re_yjp17); end else begin $fwrite(tri_report, "Item17 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per17, gol_re_yjp17, dut_re_yjp17); end end
if(col_index>=17) begin if(err_im_per17 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item17 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per17, gol_im_yjp17, dut_im_yjp17); end else begin $fwrite(tri_report, "Item17 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per17, gol_im_yjp17, dut_im_yjp17); end end

if(col_index>=18) begin if(err_re_per18 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item18 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per18, gol_re_yjp18, dut_re_yjp18); end else begin $fwrite(tri_report, "Item18 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per18, gol_re_yjp18, dut_re_yjp18); end end
if(col_index>=18) begin if(err_im_per18 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item18 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per18, gol_im_yjp18, dut_im_yjp18); end else begin $fwrite(tri_report, "Item18 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per18, gol_im_yjp18, dut_im_yjp18); end end

if(col_index>=19) begin if(err_re_per19 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item19 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per19, gol_re_yjp19, dut_re_yjp19); end else begin $fwrite(tri_report, "Item19 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per19, gol_re_yjp19, dut_re_yjp19); end end
if(col_index>=19) begin if(err_im_per19 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item19 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per19, gol_im_yjp19, dut_im_yjp19); end else begin $fwrite(tri_report, "Item19 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per19, gol_im_yjp19, dut_im_yjp19); end end

if(col_index>=20) begin if(err_re_per20 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item20 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per20, gol_re_yjp20, dut_re_yjp20); end else begin $fwrite(tri_report, "Item20 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per20, gol_re_yjp20, dut_re_yjp20); end end
if(col_index>=20) begin if(err_im_per20 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item20 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per20, gol_im_yjp20, dut_im_yjp20); end else begin $fwrite(tri_report, "Item20 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per20, gol_im_yjp20, dut_im_yjp20); end end

if(col_index>=21) begin if(err_re_per21 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item21 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per21, gol_re_yjp21, dut_re_yjp21); end else begin $fwrite(tri_report, "Item21 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per21, gol_re_yjp21, dut_re_yjp21); end end
if(col_index>=21) begin if(err_im_per21 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item21 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per21, gol_im_yjp21, dut_im_yjp21); end else begin $fwrite(tri_report, "Item21 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per21, gol_im_yjp21, dut_im_yjp21); end end

if(col_index>=22) begin if(err_re_per22 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item22 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per22, gol_re_yjp22, dut_re_yjp22); end else begin $fwrite(tri_report, "Item22 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per22, gol_re_yjp22, dut_re_yjp22); end end
if(col_index>=22) begin if(err_im_per22 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item22 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per22, gol_im_yjp22, dut_im_yjp22); end else begin $fwrite(tri_report, "Item22 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per22, gol_im_yjp22, dut_im_yjp22); end end

if(col_index>=23) begin if(err_re_per23 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item23 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per23, gol_re_yjp23, dut_re_yjp23); end else begin $fwrite(tri_report, "Item23 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per23, gol_re_yjp23, dut_re_yjp23); end end
if(col_index>=23) begin if(err_im_per23 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item23 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per23, gol_im_yjp23, dut_im_yjp23); end else begin $fwrite(tri_report, "Item23 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per23, gol_im_yjp23, dut_im_yjp23); end end

if(col_index>=24) begin if(err_re_per24 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item24 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per24, gol_re_yjp24, dut_re_yjp24); end else begin $fwrite(tri_report, "Item24 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per24, gol_re_yjp24, dut_re_yjp24); end end
if(col_index>=24) begin if(err_im_per24 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item24 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per24, gol_im_yjp24, dut_im_yjp24); end else begin $fwrite(tri_report, "Item24 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per24, gol_im_yjp24, dut_im_yjp24); end end

if(col_index>=25) begin if(err_re_per25 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item25 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per25, gol_re_yjp25, dut_re_yjp25); end else begin $fwrite(tri_report, "Item25 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per25, gol_re_yjp25, dut_re_yjp25); end end
if(col_index>=25) begin if(err_im_per25 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item25 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per25, gol_im_yjp25, dut_im_yjp25); end else begin $fwrite(tri_report, "Item25 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per25, gol_im_yjp25, dut_im_yjp25); end end

if(col_index>=26) begin if(err_re_per26 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item26 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per26, gol_re_yjp26, dut_re_yjp26); end else begin $fwrite(tri_report, "Item26 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per26, gol_re_yjp26, dut_re_yjp26); end end
if(col_index>=26) begin if(err_im_per26 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item26 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per26, gol_im_yjp26, dut_im_yjp26); end else begin $fwrite(tri_report, "Item26 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per26, gol_im_yjp26, dut_im_yjp26); end end

if(col_index>=27) begin if(err_re_per27 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item27 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per27, gol_re_yjp27, dut_re_yjp27); end else begin $fwrite(tri_report, "Item27 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per27, gol_re_yjp27, dut_re_yjp27); end end
if(col_index>=27) begin if(err_im_per27 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item27 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per27, gol_im_yjp27, dut_im_yjp27); end else begin $fwrite(tri_report, "Item27 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per27, gol_im_yjp27, dut_im_yjp27); end end

if(col_index>=28) begin if(err_re_per28 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item28 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per28, gol_re_yjp28, dut_re_yjp28); end else begin $fwrite(tri_report, "Item28 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per28, gol_re_yjp28, dut_re_yjp28); end end
if(col_index>=28) begin if(err_im_per28 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item28 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per28, gol_im_yjp28, dut_im_yjp28); end else begin $fwrite(tri_report, "Item28 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per28, gol_im_yjp28, dut_im_yjp28); end end

if(col_index>=29) begin if(err_re_per29 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item29 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per29, gol_re_yjp29, dut_re_yjp29); end else begin $fwrite(tri_report, "Item29 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per29, gol_re_yjp29, dut_re_yjp29); end end
if(col_index>=29) begin if(err_im_per29 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item29 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per29, gol_im_yjp29, dut_im_yjp29); end else begin $fwrite(tri_report, "Item29 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per29, gol_im_yjp29, dut_im_yjp29); end end

if(col_index>=30) begin if(err_re_per30 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item30 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per30, gol_re_yjp30, dut_re_yjp30); end else begin $fwrite(tri_report, "Item30 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per30, gol_re_yjp30, dut_re_yjp30); end end
if(col_index>=30) begin if(err_im_per30 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item30 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per30, gol_im_yjp30, dut_im_yjp30); end else begin $fwrite(tri_report, "Item30 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per30, gol_im_yjp30, dut_im_yjp30); end end

if(col_index>=31) begin if(err_re_per31 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item31 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per31, gol_re_yjp31, dut_re_yjp31); end else begin $fwrite(tri_report, "Item31 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per31, gol_re_yjp31, dut_re_yjp31); end end
if(col_index>=31) begin if(err_im_per31 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item31 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per31, gol_im_yjp31, dut_im_yjp31); end else begin $fwrite(tri_report, "Item31 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per31, gol_im_yjp31, dut_im_yjp31); end end

if(col_index>=32) begin if(err_re_per32 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item32 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per32, gol_re_yjp32, dut_re_yjp32); end else begin $fwrite(tri_report, "Item32 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per32, gol_re_yjp32, dut_re_yjp32); end end
if(col_index>=32) begin if(err_im_per32 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item32 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per32, gol_im_yjp32, dut_im_yjp32); end else begin $fwrite(tri_report, "Item32 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per32, gol_im_yjp32, dut_im_yjp32); end end

if(col_index>=33) begin if(err_re_per33 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item33 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per33, gol_re_yjp33, dut_re_yjp33); end else begin $fwrite(tri_report, "Item33 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per33, gol_re_yjp33, dut_re_yjp33); end end
if(col_index>=33) begin if(err_im_per33 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item33 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per33, gol_im_yjp33, dut_im_yjp33); end else begin $fwrite(tri_report, "Item33 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per33, gol_im_yjp33, dut_im_yjp33); end end

if(col_index>=34) begin if(err_re_per34 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item34 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per34, gol_re_yjp34, dut_re_yjp34); end else begin $fwrite(tri_report, "Item34 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per34, gol_re_yjp34, dut_re_yjp34); end end
if(col_index>=34) begin if(err_im_per34 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item34 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per34, gol_im_yjp34, dut_im_yjp34); end else begin $fwrite(tri_report, "Item34 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per34, gol_im_yjp34, dut_im_yjp34); end end

if(col_index>=35) begin if(err_re_per35 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item35 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per35, gol_re_yjp35, dut_re_yjp35); end else begin $fwrite(tri_report, "Item35 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per35, gol_re_yjp35, dut_re_yjp35); end end
if(col_index>=35) begin if(err_im_per35 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item35 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per35, gol_im_yjp35, dut_im_yjp35); end else begin $fwrite(tri_report, "Item35 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per35, gol_im_yjp35, dut_im_yjp35); end end

if(col_index>=36) begin if(err_re_per36 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item36 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per36, gol_re_yjp36, dut_re_yjp36); end else begin $fwrite(tri_report, "Item36 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per36, gol_re_yjp36, dut_re_yjp36); end end
if(col_index>=36) begin if(err_im_per36 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item36 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per36, gol_im_yjp36, dut_im_yjp36); end else begin $fwrite(tri_report, "Item36 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per36, gol_im_yjp36, dut_im_yjp36); end end

if(col_index>=37) begin if(err_re_per37 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item37 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per37, gol_re_yjp37, dut_re_yjp37); end else begin $fwrite(tri_report, "Item37 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per37, gol_re_yjp37, dut_re_yjp37); end end
if(col_index>=37) begin if(err_im_per37 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item37 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per37, gol_im_yjp37, dut_im_yjp37); end else begin $fwrite(tri_report, "Item37 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per37, gol_im_yjp37, dut_im_yjp37); end end

if(col_index>=38) begin if(err_re_per38 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item38 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per38, gol_re_yjp38, dut_re_yjp38); end else begin $fwrite(tri_report, "Item38 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per38, gol_re_yjp38, dut_re_yjp38); end end
if(col_index>=38) begin if(err_im_per38 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item38 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per38, gol_im_yjp38, dut_im_yjp38); end else begin $fwrite(tri_report, "Item38 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per38, gol_im_yjp38, dut_im_yjp38); end end

if(col_index>=39) begin if(err_re_per39 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item39 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per39, gol_re_yjp39, dut_re_yjp39); end else begin $fwrite(tri_report, "Item39 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per39, gol_re_yjp39, dut_re_yjp39); end end
if(col_index>=39) begin if(err_im_per39 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item39 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per39, gol_im_yjp39, dut_im_yjp39); end else begin $fwrite(tri_report, "Item39 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per39, gol_im_yjp39, dut_im_yjp39); end end

if(col_index>=40) begin if(err_re_per40 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item40 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per40, gol_re_yjp40, dut_re_yjp40); end else begin $fwrite(tri_report, "Item40 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per40, gol_re_yjp40, dut_re_yjp40); end end
if(col_index>=40) begin if(err_im_per40 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item40 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per40, gol_im_yjp40, dut_im_yjp40); end else begin $fwrite(tri_report, "Item40 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per40, gol_im_yjp40, dut_im_yjp40); end end

if(col_index>=41) begin if(err_re_per41 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item41 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per41, gol_re_yjp41, dut_re_yjp41); end else begin $fwrite(tri_report, "Item41 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per41, gol_re_yjp41, dut_re_yjp41); end end
if(col_index>=41) begin if(err_im_per41 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item41 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per41, gol_im_yjp41, dut_im_yjp41); end else begin $fwrite(tri_report, "Item41 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per41, gol_im_yjp41, dut_im_yjp41); end end

if(col_index>=42) begin if(err_re_per42 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item42 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per42, gol_re_yjp42, dut_re_yjp42); end else begin $fwrite(tri_report, "Item42 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per42, gol_re_yjp42, dut_re_yjp42); end end
if(col_index>=42) begin if(err_im_per42 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item42 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per42, gol_im_yjp42, dut_im_yjp42); end else begin $fwrite(tri_report, "Item42 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per42, gol_im_yjp42, dut_im_yjp42); end end

if(col_index>=43) begin if(err_re_per43 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item43 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per43, gol_re_yjp43, dut_re_yjp43); end else begin $fwrite(tri_report, "Item43 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per43, gol_re_yjp43, dut_re_yjp43); end end
if(col_index>=43) begin if(err_im_per43 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item43 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per43, gol_im_yjp43, dut_im_yjp43); end else begin $fwrite(tri_report, "Item43 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per43, gol_im_yjp43, dut_im_yjp43); end end

if(col_index>=44) begin if(err_re_per44 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item44 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per44, gol_re_yjp44, dut_re_yjp44); end else begin $fwrite(tri_report, "Item44 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per44, gol_re_yjp44, dut_re_yjp44); end end
if(col_index>=44) begin if(err_im_per44 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item44 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per44, gol_im_yjp44, dut_im_yjp44); end else begin $fwrite(tri_report, "Item44 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per44, gol_im_yjp44, dut_im_yjp44); end end

if(col_index>=45) begin if(err_re_per45 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item45 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per45, gol_re_yjp45, dut_re_yjp45); end else begin $fwrite(tri_report, "Item45 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per45, gol_re_yjp45, dut_re_yjp45); end end
if(col_index>=45) begin if(err_im_per45 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item45 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per45, gol_im_yjp45, dut_im_yjp45); end else begin $fwrite(tri_report, "Item45 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per45, gol_im_yjp45, dut_im_yjp45); end end

if(col_index>=46) begin if(err_re_per46 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item46 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per46, gol_re_yjp46, dut_re_yjp46); end else begin $fwrite(tri_report, "Item46 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per46, gol_re_yjp46, dut_re_yjp46); end end
if(col_index>=46) begin if(err_im_per46 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item46 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per46, gol_im_yjp46, dut_im_yjp46); end else begin $fwrite(tri_report, "Item46 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per46, gol_im_yjp46, dut_im_yjp46); end end

if(col_index>=47) begin if(err_re_per47 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item47 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per47, gol_re_yjp47, dut_re_yjp47); end else begin $fwrite(tri_report, "Item47 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per47, gol_re_yjp47, dut_re_yjp47); end end
if(col_index>=47) begin if(err_im_per47 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item47 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per47, gol_im_yjp47, dut_im_yjp47); end else begin $fwrite(tri_report, "Item47 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per47, gol_im_yjp47, dut_im_yjp47); end end

if(col_index>=48) begin if(err_re_per48 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item48 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per48, gol_re_yjp48, dut_re_yjp48); end else begin $fwrite(tri_report, "Item48 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per48, gol_re_yjp48, dut_re_yjp48); end end
if(col_index>=48) begin if(err_im_per48 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item48 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per48, gol_im_yjp48, dut_im_yjp48); end else begin $fwrite(tri_report, "Item48 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per48, gol_im_yjp48, dut_im_yjp48); end end

if(col_index>=49) begin if(err_re_per49 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item49 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per49, gol_re_yjp49, dut_re_yjp49); end else begin $fwrite(tri_report, "Item49 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per49, gol_re_yjp49, dut_re_yjp49); end end
if(col_index>=49) begin if(err_im_per49 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item49 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per49, gol_im_yjp49, dut_im_yjp49); end else begin $fwrite(tri_report, "Item49 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per49, gol_im_yjp49, dut_im_yjp49); end end

if(col_index>=50) begin if(err_re_per50 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item50 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per50, gol_re_yjp50, dut_re_yjp50); end else begin $fwrite(tri_report, "Item50 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per50, gol_re_yjp50, dut_re_yjp50); end end
if(col_index>=50) begin if(err_im_per50 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item50 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per50, gol_im_yjp50, dut_im_yjp50); end else begin $fwrite(tri_report, "Item50 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per50, gol_im_yjp50, dut_im_yjp50); end end

if(col_index>=51) begin if(err_re_per51 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item51 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per51, gol_re_yjp51, dut_re_yjp51); end else begin $fwrite(tri_report, "Item51 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per51, gol_re_yjp51, dut_re_yjp51); end end
if(col_index>=51) begin if(err_im_per51 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item51 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per51, gol_im_yjp51, dut_im_yjp51); end else begin $fwrite(tri_report, "Item51 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per51, gol_im_yjp51, dut_im_yjp51); end end

if(col_index>=52) begin if(err_re_per52 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item52 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per52, gol_re_yjp52, dut_re_yjp52); end else begin $fwrite(tri_report, "Item52 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per52, gol_re_yjp52, dut_re_yjp52); end end
if(col_index>=52) begin if(err_im_per52 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item52 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per52, gol_im_yjp52, dut_im_yjp52); end else begin $fwrite(tri_report, "Item52 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per52, gol_im_yjp52, dut_im_yjp52); end end

if(col_index>=53) begin if(err_re_per53 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item53 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per53, gol_re_yjp53, dut_re_yjp53); end else begin $fwrite(tri_report, "Item53 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per53, gol_re_yjp53, dut_re_yjp53); end end
if(col_index>=53) begin if(err_im_per53 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item53 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per53, gol_im_yjp53, dut_im_yjp53); end else begin $fwrite(tri_report, "Item53 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per53, gol_im_yjp53, dut_im_yjp53); end end

if(col_index>=54) begin if(err_re_per54 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item54 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per54, gol_re_yjp54, dut_re_yjp54); end else begin $fwrite(tri_report, "Item54 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per54, gol_re_yjp54, dut_re_yjp54); end end
if(col_index>=54) begin if(err_im_per54 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item54 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per54, gol_im_yjp54, dut_im_yjp54); end else begin $fwrite(tri_report, "Item54 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per54, gol_im_yjp54, dut_im_yjp54); end end

if(col_index>=55) begin if(err_re_per55 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item55 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per55, gol_re_yjp55, dut_re_yjp55); end else begin $fwrite(tri_report, "Item55 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per55, gol_re_yjp55, dut_re_yjp55); end end
if(col_index>=55) begin if(err_im_per55 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item55 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per55, gol_im_yjp55, dut_im_yjp55); end else begin $fwrite(tri_report, "Item55 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per55, gol_im_yjp55, dut_im_yjp55); end end

if(col_index>=56) begin if(err_re_per56 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item56 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per56, gol_re_yjp56, dut_re_yjp56); end else begin $fwrite(tri_report, "Item56 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per56, gol_re_yjp56, dut_re_yjp56); end end
if(col_index>=56) begin if(err_im_per56 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item56 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per56, gol_im_yjp56, dut_im_yjp56); end else begin $fwrite(tri_report, "Item56 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per56, gol_im_yjp56, dut_im_yjp56); end end

if(col_index>=57) begin if(err_re_per57 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item57 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per57, gol_re_yjp57, dut_re_yjp57); end else begin $fwrite(tri_report, "Item57 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per57, gol_re_yjp57, dut_re_yjp57); end end
if(col_index>=57) begin if(err_im_per57 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item57 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per57, gol_im_yjp57, dut_im_yjp57); end else begin $fwrite(tri_report, "Item57 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per57, gol_im_yjp57, dut_im_yjp57); end end

if(col_index>=58) begin if(err_re_per58 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item58 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per58, gol_re_yjp58, dut_re_yjp58); end else begin $fwrite(tri_report, "Item58 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per58, gol_re_yjp58, dut_re_yjp58); end end
if(col_index>=58) begin if(err_im_per58 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item58 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per58, gol_im_yjp58, dut_im_yjp58); end else begin $fwrite(tri_report, "Item58 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per58, gol_im_yjp58, dut_im_yjp58); end end

if(col_index>=59) begin if(err_re_per59 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item59 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per59, gol_re_yjp59, dut_re_yjp59); end else begin $fwrite(tri_report, "Item59 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per59, gol_re_yjp59, dut_re_yjp59); end end
if(col_index>=59) begin if(err_im_per59 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item59 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per59, gol_im_yjp59, dut_im_yjp59); end else begin $fwrite(tri_report, "Item59 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per59, gol_im_yjp59, dut_im_yjp59); end end

if(col_index>=60) begin if(err_re_per60 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item60 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per60, gol_re_yjp60, dut_re_yjp60); end else begin $fwrite(tri_report, "Item60 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per60, gol_re_yjp60, dut_re_yjp60); end end
if(col_index>=60) begin if(err_im_per60 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item60 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per60, gol_im_yjp60, dut_im_yjp60); end else begin $fwrite(tri_report, "Item60 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per60, gol_im_yjp60, dut_im_yjp60); end end

if(col_index>=61) begin if(err_re_per61 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item61 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per61, gol_re_yjp61, dut_re_yjp61); end else begin $fwrite(tri_report, "Item61 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per61, gol_re_yjp61, dut_re_yjp61); end end
if(col_index>=61) begin if(err_im_per61 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item61 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per61, gol_im_yjp61, dut_im_yjp61); end else begin $fwrite(tri_report, "Item61 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per61, gol_im_yjp61, dut_im_yjp61); end end

if(col_index>=62) begin if(err_re_per62 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item62 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per62, gol_re_yjp62, dut_re_yjp62); end else begin $fwrite(tri_report, "Item62 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per62, gol_re_yjp62, dut_re_yjp62); end end
if(col_index>=62) begin if(err_im_per62 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item62 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per62, gol_im_yjp62, dut_im_yjp62); end else begin $fwrite(tri_report, "Item62 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per62, gol_im_yjp62, dut_im_yjp62); end end

if(col_index>=63) begin if(err_re_per63 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item63 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per63, gol_re_yjp63, dut_re_yjp63); end else begin $fwrite(tri_report, "Item63 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per63, gol_re_yjp63, dut_re_yjp63); end end
if(col_index>=63) begin if(err_im_per63 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item63 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per63, gol_im_yjp63, dut_im_yjp63); end else begin $fwrite(tri_report, "Item63 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per63, gol_im_yjp63, dut_im_yjp63); end end

if(col_index>=64) begin if(err_re_per64 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item64 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per64, gol_re_yjp64, dut_re_yjp64); end else begin $fwrite(tri_report, "Item64 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per64, gol_re_yjp64, dut_re_yjp64); end end
if(col_index>=64) begin if(err_im_per64 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item64 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per64, gol_im_yjp64, dut_im_yjp64); end else begin $fwrite(tri_report, "Item64 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per64, gol_im_yjp64, dut_im_yjp64); end end

if(col_index>=65) begin if(err_re_per65 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item65 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per65, gol_re_yjp65, dut_re_yjp65); end else begin $fwrite(tri_report, "Item65 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per65, gol_re_yjp65, dut_re_yjp65); end end
if(col_index>=65) begin if(err_im_per65 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item65 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per65, gol_im_yjp65, dut_im_yjp65); end else begin $fwrite(tri_report, "Item65 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per65, gol_im_yjp65, dut_im_yjp65); end end

if(col_index>=66) begin if(err_re_per66 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item66 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per66, gol_re_yjp66, dut_re_yjp66); end else begin $fwrite(tri_report, "Item66 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per66, gol_re_yjp66, dut_re_yjp66); end end
if(col_index>=66) begin if(err_im_per66 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item66 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per66, gol_im_yjp66, dut_im_yjp66); end else begin $fwrite(tri_report, "Item66 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per66, gol_im_yjp66, dut_im_yjp66); end end

if(col_index>=67) begin if(err_re_per67 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item67 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per67, gol_re_yjp67, dut_re_yjp67); end else begin $fwrite(tri_report, "Item67 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per67, gol_re_yjp67, dut_re_yjp67); end end
if(col_index>=67) begin if(err_im_per67 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item67 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per67, gol_im_yjp67, dut_im_yjp67); end else begin $fwrite(tri_report, "Item67 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per67, gol_im_yjp67, dut_im_yjp67); end end

if(col_index>=68) begin if(err_re_per68 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item68 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per68, gol_re_yjp68, dut_re_yjp68); end else begin $fwrite(tri_report, "Item68 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per68, gol_re_yjp68, dut_re_yjp68); end end
if(col_index>=68) begin if(err_im_per68 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item68 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per68, gol_im_yjp68, dut_im_yjp68); end else begin $fwrite(tri_report, "Item68 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per68, gol_im_yjp68, dut_im_yjp68); end end

if(col_index>=69) begin if(err_re_per69 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item69 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per69, gol_re_yjp69, dut_re_yjp69); end else begin $fwrite(tri_report, "Item69 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per69, gol_re_yjp69, dut_re_yjp69); end end
if(col_index>=69) begin if(err_im_per69 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item69 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per69, gol_im_yjp69, dut_im_yjp69); end else begin $fwrite(tri_report, "Item69 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per69, gol_im_yjp69, dut_im_yjp69); end end

if(col_index>=70) begin if(err_re_per70 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item70 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per70, gol_re_yjp70, dut_re_yjp70); end else begin $fwrite(tri_report, "Item70 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per70, gol_re_yjp70, dut_re_yjp70); end end
if(col_index>=70) begin if(err_im_per70 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item70 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per70, gol_im_yjp70, dut_im_yjp70); end else begin $fwrite(tri_report, "Item70 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per70, gol_im_yjp70, dut_im_yjp70); end end

if(col_index>=71) begin if(err_re_per71 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item71 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per71, gol_re_yjp71, dut_re_yjp71); end else begin $fwrite(tri_report, "Item71 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per71, gol_re_yjp71, dut_re_yjp71); end end
if(col_index>=71) begin if(err_im_per71 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item71 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per71, gol_im_yjp71, dut_im_yjp71); end else begin $fwrite(tri_report, "Item71 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per71, gol_im_yjp71, dut_im_yjp71); end end

if(col_index>=72) begin if(err_re_per72 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item72 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per72, gol_re_yjp72, dut_re_yjp72); end else begin $fwrite(tri_report, "Item72 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per72, gol_re_yjp72, dut_re_yjp72); end end
if(col_index>=72) begin if(err_im_per72 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item72 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per72, gol_im_yjp72, dut_im_yjp72); end else begin $fwrite(tri_report, "Item72 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per72, gol_im_yjp72, dut_im_yjp72); end end

if(col_index>=73) begin if(err_re_per73 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item73 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per73, gol_re_yjp73, dut_re_yjp73); end else begin $fwrite(tri_report, "Item73 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per73, gol_re_yjp73, dut_re_yjp73); end end
if(col_index>=73) begin if(err_im_per73 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item73 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per73, gol_im_yjp73, dut_im_yjp73); end else begin $fwrite(tri_report, "Item73 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per73, gol_im_yjp73, dut_im_yjp73); end end

if(col_index>=74) begin if(err_re_per74 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item74 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per74, gol_re_yjp74, dut_re_yjp74); end else begin $fwrite(tri_report, "Item74 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per74, gol_re_yjp74, dut_re_yjp74); end end
if(col_index>=74) begin if(err_im_per74 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item74 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per74, gol_im_yjp74, dut_im_yjp74); end else begin $fwrite(tri_report, "Item74 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per74, gol_im_yjp74, dut_im_yjp74); end end

if(col_index>=75) begin if(err_re_per75 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item75 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per75, gol_re_yjp75, dut_re_yjp75); end else begin $fwrite(tri_report, "Item75 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per75, gol_re_yjp75, dut_re_yjp75); end end
if(col_index>=75) begin if(err_im_per75 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item75 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per75, gol_im_yjp75, dut_im_yjp75); end else begin $fwrite(tri_report, "Item75 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per75, gol_im_yjp75, dut_im_yjp75); end end

if(col_index>=76) begin if(err_re_per76 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item76 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per76, gol_re_yjp76, dut_re_yjp76); end else begin $fwrite(tri_report, "Item76 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per76, gol_re_yjp76, dut_re_yjp76); end end
if(col_index>=76) begin if(err_im_per76 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item76 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per76, gol_im_yjp76, dut_im_yjp76); end else begin $fwrite(tri_report, "Item76 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per76, gol_im_yjp76, dut_im_yjp76); end end

if(col_index>=77) begin if(err_re_per77 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item77 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per77, gol_re_yjp77, dut_re_yjp77); end else begin $fwrite(tri_report, "Item77 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per77, gol_re_yjp77, dut_re_yjp77); end end
if(col_index>=77) begin if(err_im_per77 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item77 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per77, gol_im_yjp77, dut_im_yjp77); end else begin $fwrite(tri_report, "Item77 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per77, gol_im_yjp77, dut_im_yjp77); end end

if(col_index>=78) begin if(err_re_per78 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item78 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per78, gol_re_yjp78, dut_re_yjp78); end else begin $fwrite(tri_report, "Item78 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per78, gol_re_yjp78, dut_re_yjp78); end end
if(col_index>=78) begin if(err_im_per78 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item78 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per78, gol_im_yjp78, dut_im_yjp78); end else begin $fwrite(tri_report, "Item78 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per78, gol_im_yjp78, dut_im_yjp78); end end

if(col_index>=79) begin if(err_re_per79 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item79 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per79, gol_re_yjp79, dut_re_yjp79); end else begin $fwrite(tri_report, "Item79 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per79, gol_re_yjp79, dut_re_yjp79); end end
if(col_index>=79) begin if(err_im_per79 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item79 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per79, gol_im_yjp79, dut_im_yjp79); end else begin $fwrite(tri_report, "Item79 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per79, gol_im_yjp79, dut_im_yjp79); end end

if(col_index>=80) begin if(err_re_per80 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item80 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per80, gol_re_yjp80, dut_re_yjp80); end else begin $fwrite(tri_report, "Item80 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per80, gol_re_yjp80, dut_re_yjp80); end end
if(col_index>=80) begin if(err_im_per80 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item80 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per80, gol_im_yjp80, dut_im_yjp80); end else begin $fwrite(tri_report, "Item80 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per80, gol_im_yjp80, dut_im_yjp80); end end

if(col_index>=81) begin if(err_re_per81 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item81 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per81, gol_re_yjp81, dut_re_yjp81); end else begin $fwrite(tri_report, "Item81 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per81, gol_re_yjp81, dut_re_yjp81); end end
if(col_index>=81) begin if(err_im_per81 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item81 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per81, gol_im_yjp81, dut_im_yjp81); end else begin $fwrite(tri_report, "Item81 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per81, gol_im_yjp81, dut_im_yjp81); end end

if(col_index>=82) begin if(err_re_per82 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item82 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per82, gol_re_yjp82, dut_re_yjp82); end else begin $fwrite(tri_report, "Item82 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per82, gol_re_yjp82, dut_re_yjp82); end end
if(col_index>=82) begin if(err_im_per82 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item82 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per82, gol_im_yjp82, dut_im_yjp82); end else begin $fwrite(tri_report, "Item82 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per82, gol_im_yjp82, dut_im_yjp82); end end

if(col_index>=83) begin if(err_re_per83 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item83 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per83, gol_re_yjp83, dut_re_yjp83); end else begin $fwrite(tri_report, "Item83 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per83, gol_re_yjp83, dut_re_yjp83); end end
if(col_index>=83) begin if(err_im_per83 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item83 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per83, gol_im_yjp83, dut_im_yjp83); end else begin $fwrite(tri_report, "Item83 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per83, gol_im_yjp83, dut_im_yjp83); end end

if(col_index>=84) begin if(err_re_per84 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item84 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per84, gol_re_yjp84, dut_re_yjp84); end else begin $fwrite(tri_report, "Item84 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per84, gol_re_yjp84, dut_re_yjp84); end end
if(col_index>=84) begin if(err_im_per84 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item84 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per84, gol_im_yjp84, dut_im_yjp84); end else begin $fwrite(tri_report, "Item84 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per84, gol_im_yjp84, dut_im_yjp84); end end

if(col_index>=85) begin if(err_re_per85 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item85 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per85, gol_re_yjp85, dut_re_yjp85); end else begin $fwrite(tri_report, "Item85 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per85, gol_re_yjp85, dut_re_yjp85); end end
if(col_index>=85) begin if(err_im_per85 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item85 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per85, gol_im_yjp85, dut_im_yjp85); end else begin $fwrite(tri_report, "Item85 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per85, gol_im_yjp85, dut_im_yjp85); end end

if(col_index>=86) begin if(err_re_per86 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item86 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per86, gol_re_yjp86, dut_re_yjp86); end else begin $fwrite(tri_report, "Item86 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per86, gol_re_yjp86, dut_re_yjp86); end end
if(col_index>=86) begin if(err_im_per86 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item86 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per86, gol_im_yjp86, dut_im_yjp86); end else begin $fwrite(tri_report, "Item86 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per86, gol_im_yjp86, dut_im_yjp86); end end

if(col_index>=87) begin if(err_re_per87 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item87 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per87, gol_re_yjp87, dut_re_yjp87); end else begin $fwrite(tri_report, "Item87 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per87, gol_re_yjp87, dut_re_yjp87); end end
if(col_index>=87) begin if(err_im_per87 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item87 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per87, gol_im_yjp87, dut_im_yjp87); end else begin $fwrite(tri_report, "Item87 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per87, gol_im_yjp87, dut_im_yjp87); end end

if(col_index>=88) begin if(err_re_per88 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item88 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per88, gol_re_yjp88, dut_re_yjp88); end else begin $fwrite(tri_report, "Item88 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per88, gol_re_yjp88, dut_re_yjp88); end end
if(col_index>=88) begin if(err_im_per88 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item88 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per88, gol_im_yjp88, dut_im_yjp88); end else begin $fwrite(tri_report, "Item88 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per88, gol_im_yjp88, dut_im_yjp88); end end

if(col_index>=89) begin if(err_re_per89 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item89 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per89, gol_re_yjp89, dut_re_yjp89); end else begin $fwrite(tri_report, "Item89 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per89, gol_re_yjp89, dut_re_yjp89); end end
if(col_index>=89) begin if(err_im_per89 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item89 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per89, gol_im_yjp89, dut_im_yjp89); end else begin $fwrite(tri_report, "Item89 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per89, gol_im_yjp89, dut_im_yjp89); end end

if(col_index>=90) begin if(err_re_per90 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item90 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per90, gol_re_yjp90, dut_re_yjp90); end else begin $fwrite(tri_report, "Item90 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per90, gol_re_yjp90, dut_re_yjp90); end end
if(col_index>=90) begin if(err_im_per90 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item90 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per90, gol_im_yjp90, dut_im_yjp90); end else begin $fwrite(tri_report, "Item90 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per90, gol_im_yjp90, dut_im_yjp90); end end

if(col_index>=91) begin if(err_re_per91 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item91 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per91, gol_re_yjp91, dut_re_yjp91); end else begin $fwrite(tri_report, "Item91 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per91, gol_re_yjp91, dut_re_yjp91); end end
if(col_index>=91) begin if(err_im_per91 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item91 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per91, gol_im_yjp91, dut_im_yjp91); end else begin $fwrite(tri_report, "Item91 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per91, gol_im_yjp91, dut_im_yjp91); end end

if(col_index>=92) begin if(err_re_per92 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item92 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per92, gol_re_yjp92, dut_re_yjp92); end else begin $fwrite(tri_report, "Item92 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per92, gol_re_yjp92, dut_re_yjp92); end end
if(col_index>=92) begin if(err_im_per92 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item92 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per92, gol_im_yjp92, dut_im_yjp92); end else begin $fwrite(tri_report, "Item92 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per92, gol_im_yjp92, dut_im_yjp92); end end

if(col_index>=93) begin if(err_re_per93 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item93 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per93, gol_re_yjp93, dut_re_yjp93); end else begin $fwrite(tri_report, "Item93 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per93, gol_re_yjp93, dut_re_yjp93); end end
if(col_index>=93) begin if(err_im_per93 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item93 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per93, gol_im_yjp93, dut_im_yjp93); end else begin $fwrite(tri_report, "Item93 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per93, gol_im_yjp93, dut_im_yjp93); end end

if(col_index>=94) begin if(err_re_per94 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item94 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per94, gol_re_yjp94, dut_re_yjp94); end else begin $fwrite(tri_report, "Item94 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per94, gol_re_yjp94, dut_re_yjp94); end end
if(col_index>=94) begin if(err_im_per94 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item94 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per94, gol_im_yjp94, dut_im_yjp94); end else begin $fwrite(tri_report, "Item94 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per94, gol_im_yjp94, dut_im_yjp94); end end

if(col_index>=95) begin if(err_re_per95 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item95 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per95, gol_re_yjp95, dut_re_yjp95); end else begin $fwrite(tri_report, "Item95 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per95, gol_re_yjp95, dut_re_yjp95); end end
if(col_index>=95) begin if(err_im_per95 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item95 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per95, gol_im_yjp95, dut_im_yjp95); end else begin $fwrite(tri_report, "Item95 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per95, gol_im_yjp95, dut_im_yjp95); end end

if(col_index>=96) begin if(err_re_per96 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item96 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per96, gol_re_yjp96, dut_re_yjp96); end else begin $fwrite(tri_report, "Item96 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per96, gol_re_yjp96, dut_re_yjp96); end end
if(col_index>=96) begin if(err_im_per96 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item96 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per96, gol_im_yjp96, dut_im_yjp96); end else begin $fwrite(tri_report, "Item96 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per96, gol_im_yjp96, dut_im_yjp96); end end

if(col_index>=97) begin if(err_re_per97 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item97 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per97, gol_re_yjp97, dut_re_yjp97); end else begin $fwrite(tri_report, "Item97 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per97, gol_re_yjp97, dut_re_yjp97); end end
if(col_index>=97) begin if(err_im_per97 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item97 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per97, gol_im_yjp97, dut_im_yjp97); end else begin $fwrite(tri_report, "Item97 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per97, gol_im_yjp97, dut_im_yjp97); end end

if(col_index>=98) begin if(err_re_per98 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item98 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per98, gol_re_yjp98, dut_re_yjp98); end else begin $fwrite(tri_report, "Item98 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per98, gol_re_yjp98, dut_re_yjp98); end end
if(col_index>=98) begin if(err_im_per98 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item98 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per98, gol_im_yjp98, dut_im_yjp98); end else begin $fwrite(tri_report, "Item98 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per98, gol_im_yjp98, dut_im_yjp98); end end

if(col_index>=99) begin if(err_re_per99 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item99 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per99, gol_re_yjp99, dut_re_yjp99); end else begin $fwrite(tri_report, "Item99 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per99, gol_re_yjp99, dut_re_yjp99); end end
if(col_index>=99) begin if(err_im_per99 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item99 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per99, gol_im_yjp99, dut_im_yjp99); end else begin $fwrite(tri_report, "Item99 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per99, gol_im_yjp99, dut_im_yjp99); end end

if(col_index>=100) begin if(err_re_per100 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item100 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per100, gol_re_yjp100, dut_re_yjp100); end else begin $fwrite(tri_report, "Item100 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per100, gol_re_yjp100, dut_re_yjp100); end end
if(col_index>=100) begin if(err_im_per100 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item100 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per100, gol_im_yjp100, dut_im_yjp100); end else begin $fwrite(tri_report, "Item100 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per100, gol_im_yjp100, dut_im_yjp100); end end

if(col_index>=101) begin if(err_re_per101 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item101 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per101, gol_re_yjp101, dut_re_yjp101); end else begin $fwrite(tri_report, "Item101 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per101, gol_re_yjp101, dut_re_yjp101); end end
if(col_index>=101) begin if(err_im_per101 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item101 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per101, gol_im_yjp101, dut_im_yjp101); end else begin $fwrite(tri_report, "Item101 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per101, gol_im_yjp101, dut_im_yjp101); end end

if(col_index>=102) begin if(err_re_per102 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item102 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per102, gol_re_yjp102, dut_re_yjp102); end else begin $fwrite(tri_report, "Item102 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per102, gol_re_yjp102, dut_re_yjp102); end end
if(col_index>=102) begin if(err_im_per102 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item102 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per102, gol_im_yjp102, dut_im_yjp102); end else begin $fwrite(tri_report, "Item102 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per102, gol_im_yjp102, dut_im_yjp102); end end

if(col_index>=103) begin if(err_re_per103 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item103 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per103, gol_re_yjp103, dut_re_yjp103); end else begin $fwrite(tri_report, "Item103 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per103, gol_re_yjp103, dut_re_yjp103); end end
if(col_index>=103) begin if(err_im_per103 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item103 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per103, gol_im_yjp103, dut_im_yjp103); end else begin $fwrite(tri_report, "Item103 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per103, gol_im_yjp103, dut_im_yjp103); end end

if(col_index>=104) begin if(err_re_per104 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item104 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per104, gol_re_yjp104, dut_re_yjp104); end else begin $fwrite(tri_report, "Item104 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per104, gol_re_yjp104, dut_re_yjp104); end end
if(col_index>=104) begin if(err_im_per104 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item104 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per104, gol_im_yjp104, dut_im_yjp104); end else begin $fwrite(tri_report, "Item104 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per104, gol_im_yjp104, dut_im_yjp104); end end

if(col_index>=105) begin if(err_re_per105 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item105 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per105, gol_re_yjp105, dut_re_yjp105); end else begin $fwrite(tri_report, "Item105 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per105, gol_re_yjp105, dut_re_yjp105); end end
if(col_index>=105) begin if(err_im_per105 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item105 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per105, gol_im_yjp105, dut_im_yjp105); end else begin $fwrite(tri_report, "Item105 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per105, gol_im_yjp105, dut_im_yjp105); end end

if(col_index>=106) begin if(err_re_per106 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item106 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per106, gol_re_yjp106, dut_re_yjp106); end else begin $fwrite(tri_report, "Item106 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per106, gol_re_yjp106, dut_re_yjp106); end end
if(col_index>=106) begin if(err_im_per106 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item106 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per106, gol_im_yjp106, dut_im_yjp106); end else begin $fwrite(tri_report, "Item106 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per106, gol_im_yjp106, dut_im_yjp106); end end

if(col_index>=107) begin if(err_re_per107 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item107 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per107, gol_re_yjp107, dut_re_yjp107); end else begin $fwrite(tri_report, "Item107 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per107, gol_re_yjp107, dut_re_yjp107); end end
if(col_index>=107) begin if(err_im_per107 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item107 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per107, gol_im_yjp107, dut_im_yjp107); end else begin $fwrite(tri_report, "Item107 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per107, gol_im_yjp107, dut_im_yjp107); end end

if(col_index>=108) begin if(err_re_per108 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item108 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per108, gol_re_yjp108, dut_re_yjp108); end else begin $fwrite(tri_report, "Item108 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per108, gol_re_yjp108, dut_re_yjp108); end end
if(col_index>=108) begin if(err_im_per108 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item108 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per108, gol_im_yjp108, dut_im_yjp108); end else begin $fwrite(tri_report, "Item108 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per108, gol_im_yjp108, dut_im_yjp108); end end

if(col_index>=109) begin if(err_re_per109 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item109 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per109, gol_re_yjp109, dut_re_yjp109); end else begin $fwrite(tri_report, "Item109 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per109, gol_re_yjp109, dut_re_yjp109); end end
if(col_index>=109) begin if(err_im_per109 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item109 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per109, gol_im_yjp109, dut_im_yjp109); end else begin $fwrite(tri_report, "Item109 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per109, gol_im_yjp109, dut_im_yjp109); end end

if(col_index>=110) begin if(err_re_per110 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item110 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per110, gol_re_yjp110, dut_re_yjp110); end else begin $fwrite(tri_report, "Item110 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per110, gol_re_yjp110, dut_re_yjp110); end end
if(col_index>=110) begin if(err_im_per110 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item110 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per110, gol_im_yjp110, dut_im_yjp110); end else begin $fwrite(tri_report, "Item110 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per110, gol_im_yjp110, dut_im_yjp110); end end

if(col_index>=111) begin if(err_re_per111 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item111 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per111, gol_re_yjp111, dut_re_yjp111); end else begin $fwrite(tri_report, "Item111 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per111, gol_re_yjp111, dut_re_yjp111); end end
if(col_index>=111) begin if(err_im_per111 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item111 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per111, gol_im_yjp111, dut_im_yjp111); end else begin $fwrite(tri_report, "Item111 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per111, gol_im_yjp111, dut_im_yjp111); end end

if(col_index>=112) begin if(err_re_per112 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item112 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per112, gol_re_yjp112, dut_re_yjp112); end else begin $fwrite(tri_report, "Item112 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per112, gol_re_yjp112, dut_re_yjp112); end end
if(col_index>=112) begin if(err_im_per112 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item112 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per112, gol_im_yjp112, dut_im_yjp112); end else begin $fwrite(tri_report, "Item112 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per112, gol_im_yjp112, dut_im_yjp112); end end

if(col_index>=113) begin if(err_re_per113 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item113 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per113, gol_re_yjp113, dut_re_yjp113); end else begin $fwrite(tri_report, "Item113 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per113, gol_re_yjp113, dut_re_yjp113); end end
if(col_index>=113) begin if(err_im_per113 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item113 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per113, gol_im_yjp113, dut_im_yjp113); end else begin $fwrite(tri_report, "Item113 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per113, gol_im_yjp113, dut_im_yjp113); end end

if(col_index>=114) begin if(err_re_per114 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item114 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per114, gol_re_yjp114, dut_re_yjp114); end else begin $fwrite(tri_report, "Item114 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per114, gol_re_yjp114, dut_re_yjp114); end end
if(col_index>=114) begin if(err_im_per114 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item114 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per114, gol_im_yjp114, dut_im_yjp114); end else begin $fwrite(tri_report, "Item114 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per114, gol_im_yjp114, dut_im_yjp114); end end

if(col_index>=115) begin if(err_re_per115 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item115 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per115, gol_re_yjp115, dut_re_yjp115); end else begin $fwrite(tri_report, "Item115 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per115, gol_re_yjp115, dut_re_yjp115); end end
if(col_index>=115) begin if(err_im_per115 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item115 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per115, gol_im_yjp115, dut_im_yjp115); end else begin $fwrite(tri_report, "Item115 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per115, gol_im_yjp115, dut_im_yjp115); end end

if(col_index>=116) begin if(err_re_per116 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item116 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per116, gol_re_yjp116, dut_re_yjp116); end else begin $fwrite(tri_report, "Item116 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per116, gol_re_yjp116, dut_re_yjp116); end end
if(col_index>=116) begin if(err_im_per116 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item116 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per116, gol_im_yjp116, dut_im_yjp116); end else begin $fwrite(tri_report, "Item116 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per116, gol_im_yjp116, dut_im_yjp116); end end

if(col_index>=117) begin if(err_re_per117 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item117 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per117, gol_re_yjp117, dut_re_yjp117); end else begin $fwrite(tri_report, "Item117 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per117, gol_re_yjp117, dut_re_yjp117); end end
if(col_index>=117) begin if(err_im_per117 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item117 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per117, gol_im_yjp117, dut_im_yjp117); end else begin $fwrite(tri_report, "Item117 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per117, gol_im_yjp117, dut_im_yjp117); end end

if(col_index>=118) begin if(err_re_per118 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item118 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per118, gol_re_yjp118, dut_re_yjp118); end else begin $fwrite(tri_report, "Item118 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per118, gol_re_yjp118, dut_re_yjp118); end end
if(col_index>=118) begin if(err_im_per118 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item118 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per118, gol_im_yjp118, dut_im_yjp118); end else begin $fwrite(tri_report, "Item118 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per118, gol_im_yjp118, dut_im_yjp118); end end

if(col_index>=119) begin if(err_re_per119 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item119 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per119, gol_re_yjp119, dut_re_yjp119); end else begin $fwrite(tri_report, "Item119 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per119, gol_re_yjp119, dut_re_yjp119); end end
if(col_index>=119) begin if(err_im_per119 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item119 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per119, gol_im_yjp119, dut_im_yjp119); end else begin $fwrite(tri_report, "Item119 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per119, gol_im_yjp119, dut_im_yjp119); end end

if(col_index>=120) begin if(err_re_per120 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item120 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per120, gol_re_yjp120, dut_re_yjp120); end else begin $fwrite(tri_report, "Item120 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per120, gol_re_yjp120, dut_re_yjp120); end end
if(col_index>=120) begin if(err_im_per120 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item120 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per120, gol_im_yjp120, dut_im_yjp120); end else begin $fwrite(tri_report, "Item120 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per120, gol_im_yjp120, dut_im_yjp120); end end

if(col_index>=121) begin if(err_re_per121 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item121 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per121, gol_re_yjp121, dut_re_yjp121); end else begin $fwrite(tri_report, "Item121 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per121, gol_re_yjp121, dut_re_yjp121); end end
if(col_index>=121) begin if(err_im_per121 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item121 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per121, gol_im_yjp121, dut_im_yjp121); end else begin $fwrite(tri_report, "Item121 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per121, gol_im_yjp121, dut_im_yjp121); end end

if(col_index>=122) begin if(err_re_per122 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item122 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per122, gol_re_yjp122, dut_re_yjp122); end else begin $fwrite(tri_report, "Item122 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per122, gol_re_yjp122, dut_re_yjp122); end end
if(col_index>=122) begin if(err_im_per122 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item122 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per122, gol_im_yjp122, dut_im_yjp122); end else begin $fwrite(tri_report, "Item122 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per122, gol_im_yjp122, dut_im_yjp122); end end

if(col_index>=123) begin if(err_re_per123 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item123 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per123, gol_re_yjp123, dut_re_yjp123); end else begin $fwrite(tri_report, "Item123 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per123, gol_re_yjp123, dut_re_yjp123); end end
if(col_index>=123) begin if(err_im_per123 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item123 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per123, gol_im_yjp123, dut_im_yjp123); end else begin $fwrite(tri_report, "Item123 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per123, gol_im_yjp123, dut_im_yjp123); end end

if(col_index>=124) begin if(err_re_per124 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item124 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per124, gol_re_yjp124, dut_re_yjp124); end else begin $fwrite(tri_report, "Item124 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per124, gol_re_yjp124, dut_re_yjp124); end end
if(col_index>=124) begin if(err_im_per124 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item124 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per124, gol_im_yjp124, dut_im_yjp124); end else begin $fwrite(tri_report, "Item124 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per124, gol_im_yjp124, dut_im_yjp124); end end

if(col_index>=125) begin if(err_re_per125 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item125 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per125, gol_re_yjp125, dut_re_yjp125); end else begin $fwrite(tri_report, "Item125 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per125, gol_re_yjp125, dut_re_yjp125); end end
if(col_index>=125) begin if(err_im_per125 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item125 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per125, gol_im_yjp125, dut_im_yjp125); end else begin $fwrite(tri_report, "Item125 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per125, gol_im_yjp125, dut_im_yjp125); end end

if(col_index>=126) begin if(err_re_per126 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item126 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per126, gol_re_yjp126, dut_re_yjp126); end else begin $fwrite(tri_report, "Item126 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per126, gol_re_yjp126, dut_re_yjp126); end end
if(col_index>=126) begin if(err_im_per126 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item126 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per126, gol_im_yjp126, dut_im_yjp126); end else begin $fwrite(tri_report, "Item126 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per126, gol_im_yjp126, dut_im_yjp126); end end

if(col_index>=127) begin if(err_re_per127 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item127 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per127, gol_re_yjp127, dut_re_yjp127); end else begin $fwrite(tri_report, "Item127 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per127, gol_re_yjp127, dut_re_yjp127); end end
if(col_index>=127) begin if(err_im_per127 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item127 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per127, gol_im_yjp127, dut_im_yjp127); end else begin $fwrite(tri_report, "Item127 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per127, gol_im_yjp127, dut_im_yjp127); end end

if(col_index>=128) begin if(err_re_per128 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item128 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per128, gol_re_yjp128, dut_re_yjp128); end else begin $fwrite(tri_report, "Item128 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per128, gol_re_yjp128, dut_re_yjp128); end end
if(col_index>=128) begin if(err_im_per128 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item128 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per128, gol_im_yjp128, dut_im_yjp128); end else begin $fwrite(tri_report, "Item128 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per128, gol_im_yjp128, dut_im_yjp128); end end

if(col_index>=129) begin if(err_re_per129 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item129 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per129, gol_re_yjp129, dut_re_yjp129); end else begin $fwrite(tri_report, "Item129 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per129, gol_re_yjp129, dut_re_yjp129); end end
if(col_index>=129) begin if(err_im_per129 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item129 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per129, gol_im_yjp129, dut_im_yjp129); end else begin $fwrite(tri_report, "Item129 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per129, gol_im_yjp129, dut_im_yjp129); end end

if(col_index>=130) begin if(err_re_per130 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item130 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per130, gol_re_yjp130, dut_re_yjp130); end else begin $fwrite(tri_report, "Item130 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per130, gol_re_yjp130, dut_re_yjp130); end end
if(col_index>=130) begin if(err_im_per130 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item130 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per130, gol_im_yjp130, dut_im_yjp130); end else begin $fwrite(tri_report, "Item130 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per130, gol_im_yjp130, dut_im_yjp130); end end

if(col_index>=131) begin if(err_re_per131 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item131 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per131, gol_re_yjp131, dut_re_yjp131); end else begin $fwrite(tri_report, "Item131 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per131, gol_re_yjp131, dut_re_yjp131); end end
if(col_index>=131) begin if(err_im_per131 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item131 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per131, gol_im_yjp131, dut_im_yjp131); end else begin $fwrite(tri_report, "Item131 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per131, gol_im_yjp131, dut_im_yjp131); end end

if(col_index>=132) begin if(err_re_per132 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item132 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per132, gol_re_yjp132, dut_re_yjp132); end else begin $fwrite(tri_report, "Item132 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per132, gol_re_yjp132, dut_re_yjp132); end end
if(col_index>=132) begin if(err_im_per132 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item132 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per132, gol_im_yjp132, dut_im_yjp132); end else begin $fwrite(tri_report, "Item132 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per132, gol_im_yjp132, dut_im_yjp132); end end

if(col_index>=133) begin if(err_re_per133 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item133 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per133, gol_re_yjp133, dut_re_yjp133); end else begin $fwrite(tri_report, "Item133 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per133, gol_re_yjp133, dut_re_yjp133); end end
if(col_index>=133) begin if(err_im_per133 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item133 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per133, gol_im_yjp133, dut_im_yjp133); end else begin $fwrite(tri_report, "Item133 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per133, gol_im_yjp133, dut_im_yjp133); end end

if(col_index>=134) begin if(err_re_per134 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item134 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per134, gol_re_yjp134, dut_re_yjp134); end else begin $fwrite(tri_report, "Item134 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per134, gol_re_yjp134, dut_re_yjp134); end end
if(col_index>=134) begin if(err_im_per134 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item134 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per134, gol_im_yjp134, dut_im_yjp134); end else begin $fwrite(tri_report, "Item134 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per134, gol_im_yjp134, dut_im_yjp134); end end

if(col_index>=135) begin if(err_re_per135 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item135 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per135, gol_re_yjp135, dut_re_yjp135); end else begin $fwrite(tri_report, "Item135 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per135, gol_re_yjp135, dut_re_yjp135); end end
if(col_index>=135) begin if(err_im_per135 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item135 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per135, gol_im_yjp135, dut_im_yjp135); end else begin $fwrite(tri_report, "Item135 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per135, gol_im_yjp135, dut_im_yjp135); end end

if(col_index>=136) begin if(err_re_per136 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item136 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per136, gol_re_yjp136, dut_re_yjp136); end else begin $fwrite(tri_report, "Item136 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per136, gol_re_yjp136, dut_re_yjp136); end end
if(col_index>=136) begin if(err_im_per136 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item136 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per136, gol_im_yjp136, dut_im_yjp136); end else begin $fwrite(tri_report, "Item136 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per136, gol_im_yjp136, dut_im_yjp136); end end

if(col_index>=137) begin if(err_re_per137 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item137 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per137, gol_re_yjp137, dut_re_yjp137); end else begin $fwrite(tri_report, "Item137 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per137, gol_re_yjp137, dut_re_yjp137); end end
if(col_index>=137) begin if(err_im_per137 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item137 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per137, gol_im_yjp137, dut_im_yjp137); end else begin $fwrite(tri_report, "Item137 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per137, gol_im_yjp137, dut_im_yjp137); end end

if(col_index>=138) begin if(err_re_per138 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item138 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per138, gol_re_yjp138, dut_re_yjp138); end else begin $fwrite(tri_report, "Item138 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per138, gol_re_yjp138, dut_re_yjp138); end end
if(col_index>=138) begin if(err_im_per138 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item138 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per138, gol_im_yjp138, dut_im_yjp138); end else begin $fwrite(tri_report, "Item138 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per138, gol_im_yjp138, dut_im_yjp138); end end

if(col_index>=139) begin if(err_re_per139 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item139 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per139, gol_re_yjp139, dut_re_yjp139); end else begin $fwrite(tri_report, "Item139 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per139, gol_re_yjp139, dut_re_yjp139); end end
if(col_index>=139) begin if(err_im_per139 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item139 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per139, gol_im_yjp139, dut_im_yjp139); end else begin $fwrite(tri_report, "Item139 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per139, gol_im_yjp139, dut_im_yjp139); end end

if(col_index>=140) begin if(err_re_per140 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item140 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per140, gol_re_yjp140, dut_re_yjp140); end else begin $fwrite(tri_report, "Item140 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per140, gol_re_yjp140, dut_re_yjp140); end end
if(col_index>=140) begin if(err_im_per140 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item140 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per140, gol_im_yjp140, dut_im_yjp140); end else begin $fwrite(tri_report, "Item140 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per140, gol_im_yjp140, dut_im_yjp140); end end

if(col_index>=141) begin if(err_re_per141 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item141 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per141, gol_re_yjp141, dut_re_yjp141); end else begin $fwrite(tri_report, "Item141 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per141, gol_re_yjp141, dut_re_yjp141); end end
if(col_index>=141) begin if(err_im_per141 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item141 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per141, gol_im_yjp141, dut_im_yjp141); end else begin $fwrite(tri_report, "Item141 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per141, gol_im_yjp141, dut_im_yjp141); end end

if(col_index>=142) begin if(err_re_per142 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item142 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per142, gol_re_yjp142, dut_re_yjp142); end else begin $fwrite(tri_report, "Item142 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per142, gol_re_yjp142, dut_re_yjp142); end end
if(col_index>=142) begin if(err_im_per142 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item142 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per142, gol_im_yjp142, dut_im_yjp142); end else begin $fwrite(tri_report, "Item142 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per142, gol_im_yjp142, dut_im_yjp142); end end

if(col_index>=143) begin if(err_re_per143 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item143 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per143, gol_re_yjp143, dut_re_yjp143); end else begin $fwrite(tri_report, "Item143 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per143, gol_re_yjp143, dut_re_yjp143); end end
if(col_index>=143) begin if(err_im_per143 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item143 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per143, gol_im_yjp143, dut_im_yjp143); end else begin $fwrite(tri_report, "Item143 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per143, gol_im_yjp143, dut_im_yjp143); end end

if(col_index>=144) begin if(err_re_per144 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item144 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per144, gol_re_yjp144, dut_re_yjp144); end else begin $fwrite(tri_report, "Item144 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per144, gol_re_yjp144, dut_re_yjp144); end end
if(col_index>=144) begin if(err_im_per144 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item144 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per144, gol_im_yjp144, dut_im_yjp144); end else begin $fwrite(tri_report, "Item144 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per144, gol_im_yjp144, dut_im_yjp144); end end

if(col_index>=145) begin if(err_re_per145 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item145 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per145, gol_re_yjp145, dut_re_yjp145); end else begin $fwrite(tri_report, "Item145 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per145, gol_re_yjp145, dut_re_yjp145); end end
if(col_index>=145) begin if(err_im_per145 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item145 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per145, gol_im_yjp145, dut_im_yjp145); end else begin $fwrite(tri_report, "Item145 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per145, gol_im_yjp145, dut_im_yjp145); end end

if(col_index>=146) begin if(err_re_per146 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item146 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per146, gol_re_yjp146, dut_re_yjp146); end else begin $fwrite(tri_report, "Item146 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per146, gol_re_yjp146, dut_re_yjp146); end end
if(col_index>=146) begin if(err_im_per146 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item146 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per146, gol_im_yjp146, dut_im_yjp146); end else begin $fwrite(tri_report, "Item146 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per146, gol_im_yjp146, dut_im_yjp146); end end

if(col_index>=147) begin if(err_re_per147 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item147 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per147, gol_re_yjp147, dut_re_yjp147); end else begin $fwrite(tri_report, "Item147 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per147, gol_re_yjp147, dut_re_yjp147); end end
if(col_index>=147) begin if(err_im_per147 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item147 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per147, gol_im_yjp147, dut_im_yjp147); end else begin $fwrite(tri_report, "Item147 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per147, gol_im_yjp147, dut_im_yjp147); end end

if(col_index>=148) begin if(err_re_per148 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item148 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per148, gol_re_yjp148, dut_re_yjp148); end else begin $fwrite(tri_report, "Item148 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per148, gol_re_yjp148, dut_re_yjp148); end end
if(col_index>=148) begin if(err_im_per148 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item148 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per148, gol_im_yjp148, dut_im_yjp148); end else begin $fwrite(tri_report, "Item148 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per148, gol_im_yjp148, dut_im_yjp148); end end

if(col_index>=149) begin if(err_re_per149 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item149 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per149, gol_re_yjp149, dut_re_yjp149); end else begin $fwrite(tri_report, "Item149 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per149, gol_re_yjp149, dut_re_yjp149); end end
if(col_index>=149) begin if(err_im_per149 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item149 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per149, gol_im_yjp149, dut_im_yjp149); end else begin $fwrite(tri_report, "Item149 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per149, gol_im_yjp149, dut_im_yjp149); end end

if(col_index>=150) begin if(err_re_per150 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item150 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per150, gol_re_yjp150, dut_re_yjp150); end else begin $fwrite(tri_report, "Item150 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per150, gol_re_yjp150, dut_re_yjp150); end end
if(col_index>=150) begin if(err_im_per150 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item150 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per150, gol_im_yjp150, dut_im_yjp150); end else begin $fwrite(tri_report, "Item150 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per150, gol_im_yjp150, dut_im_yjp150); end end

if(col_index>=151) begin if(err_re_per151 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item151 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per151, gol_re_yjp151, dut_re_yjp151); end else begin $fwrite(tri_report, "Item151 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per151, gol_re_yjp151, dut_re_yjp151); end end
if(col_index>=151) begin if(err_im_per151 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item151 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per151, gol_im_yjp151, dut_im_yjp151); end else begin $fwrite(tri_report, "Item151 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per151, gol_im_yjp151, dut_im_yjp151); end end

if(col_index>=152) begin if(err_re_per152 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item152 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per152, gol_re_yjp152, dut_re_yjp152); end else begin $fwrite(tri_report, "Item152 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per152, gol_re_yjp152, dut_re_yjp152); end end
if(col_index>=152) begin if(err_im_per152 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item152 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per152, gol_im_yjp152, dut_im_yjp152); end else begin $fwrite(tri_report, "Item152 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per152, gol_im_yjp152, dut_im_yjp152); end end

if(col_index>=153) begin if(err_re_per153 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item153 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per153, gol_re_yjp153, dut_re_yjp153); end else begin $fwrite(tri_report, "Item153 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per153, gol_re_yjp153, dut_re_yjp153); end end
if(col_index>=153) begin if(err_im_per153 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item153 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per153, gol_im_yjp153, dut_im_yjp153); end else begin $fwrite(tri_report, "Item153 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per153, gol_im_yjp153, dut_im_yjp153); end end

if(col_index>=154) begin if(err_re_per154 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item154 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per154, gol_re_yjp154, dut_re_yjp154); end else begin $fwrite(tri_report, "Item154 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per154, gol_re_yjp154, dut_re_yjp154); end end
if(col_index>=154) begin if(err_im_per154 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item154 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per154, gol_im_yjp154, dut_im_yjp154); end else begin $fwrite(tri_report, "Item154 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per154, gol_im_yjp154, dut_im_yjp154); end end

if(col_index>=155) begin if(err_re_per155 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item155 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per155, gol_re_yjp155, dut_re_yjp155); end else begin $fwrite(tri_report, "Item155 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per155, gol_re_yjp155, dut_re_yjp155); end end
if(col_index>=155) begin if(err_im_per155 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item155 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per155, gol_im_yjp155, dut_im_yjp155); end else begin $fwrite(tri_report, "Item155 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per155, gol_im_yjp155, dut_im_yjp155); end end

if(col_index>=156) begin if(err_re_per156 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item156 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per156, gol_re_yjp156, dut_re_yjp156); end else begin $fwrite(tri_report, "Item156 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per156, gol_re_yjp156, dut_re_yjp156); end end
if(col_index>=156) begin if(err_im_per156 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item156 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per156, gol_im_yjp156, dut_im_yjp156); end else begin $fwrite(tri_report, "Item156 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per156, gol_im_yjp156, dut_im_yjp156); end end

if(col_index>=157) begin if(err_re_per157 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item157 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per157, gol_re_yjp157, dut_re_yjp157); end else begin $fwrite(tri_report, "Item157 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per157, gol_re_yjp157, dut_re_yjp157); end end
if(col_index>=157) begin if(err_im_per157 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item157 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per157, gol_im_yjp157, dut_im_yjp157); end else begin $fwrite(tri_report, "Item157 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per157, gol_im_yjp157, dut_im_yjp157); end end

if(col_index>=158) begin if(err_re_per158 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item158 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per158, gol_re_yjp158, dut_re_yjp158); end else begin $fwrite(tri_report, "Item158 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per158, gol_re_yjp158, dut_re_yjp158); end end
if(col_index>=158) begin if(err_im_per158 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item158 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per158, gol_im_yjp158, dut_im_yjp158); end else begin $fwrite(tri_report, "Item158 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per158, gol_im_yjp158, dut_im_yjp158); end end

if(col_index>=159) begin if(err_re_per159 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item159 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per159, gol_re_yjp159, dut_re_yjp159); end else begin $fwrite(tri_report, "Item159 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per159, gol_re_yjp159, dut_re_yjp159); end end
if(col_index>=159) begin if(err_im_per159 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item159 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per159, gol_im_yjp159, dut_im_yjp159); end else begin $fwrite(tri_report, "Item159 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per159, gol_im_yjp159, dut_im_yjp159); end end

if(col_index>=160) begin if(err_re_per160 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item160 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per160, gol_re_yjp160, dut_re_yjp160); end else begin $fwrite(tri_report, "Item160 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per160, gol_re_yjp160, dut_re_yjp160); end end
if(col_index>=160) begin if(err_im_per160 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item160 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per160, gol_im_yjp160, dut_im_yjp160); end else begin $fwrite(tri_report, "Item160 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per160, gol_im_yjp160, dut_im_yjp160); end end

if(col_index>=161) begin if(err_re_per161 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item161 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per161, gol_re_yjp161, dut_re_yjp161); end else begin $fwrite(tri_report, "Item161 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per161, gol_re_yjp161, dut_re_yjp161); end end
if(col_index>=161) begin if(err_im_per161 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item161 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per161, gol_im_yjp161, dut_im_yjp161); end else begin $fwrite(tri_report, "Item161 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per161, gol_im_yjp161, dut_im_yjp161); end end

if(col_index>=162) begin if(err_re_per162 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item162 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per162, gol_re_yjp162, dut_re_yjp162); end else begin $fwrite(tri_report, "Item162 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per162, gol_re_yjp162, dut_re_yjp162); end end
if(col_index>=162) begin if(err_im_per162 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item162 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per162, gol_im_yjp162, dut_im_yjp162); end else begin $fwrite(tri_report, "Item162 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per162, gol_im_yjp162, dut_im_yjp162); end end

if(col_index>=163) begin if(err_re_per163 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item163 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per163, gol_re_yjp163, dut_re_yjp163); end else begin $fwrite(tri_report, "Item163 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per163, gol_re_yjp163, dut_re_yjp163); end end
if(col_index>=163) begin if(err_im_per163 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item163 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per163, gol_im_yjp163, dut_im_yjp163); end else begin $fwrite(tri_report, "Item163 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per163, gol_im_yjp163, dut_im_yjp163); end end

if(col_index>=164) begin if(err_re_per164 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item164 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per164, gol_re_yjp164, dut_re_yjp164); end else begin $fwrite(tri_report, "Item164 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per164, gol_re_yjp164, dut_re_yjp164); end end
if(col_index>=164) begin if(err_im_per164 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item164 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per164, gol_im_yjp164, dut_im_yjp164); end else begin $fwrite(tri_report, "Item164 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per164, gol_im_yjp164, dut_im_yjp164); end end

if(col_index>=165) begin if(err_re_per165 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item165 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per165, gol_re_yjp165, dut_re_yjp165); end else begin $fwrite(tri_report, "Item165 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per165, gol_re_yjp165, dut_re_yjp165); end end
if(col_index>=165) begin if(err_im_per165 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item165 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per165, gol_im_yjp165, dut_im_yjp165); end else begin $fwrite(tri_report, "Item165 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per165, gol_im_yjp165, dut_im_yjp165); end end

if(col_index>=166) begin if(err_re_per166 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item166 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per166, gol_re_yjp166, dut_re_yjp166); end else begin $fwrite(tri_report, "Item166 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per166, gol_re_yjp166, dut_re_yjp166); end end
if(col_index>=166) begin if(err_im_per166 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item166 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per166, gol_im_yjp166, dut_im_yjp166); end else begin $fwrite(tri_report, "Item166 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per166, gol_im_yjp166, dut_im_yjp166); end end

if(col_index>=167) begin if(err_re_per167 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item167 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per167, gol_re_yjp167, dut_re_yjp167); end else begin $fwrite(tri_report, "Item167 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per167, gol_re_yjp167, dut_re_yjp167); end end
if(col_index>=167) begin if(err_im_per167 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item167 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per167, gol_im_yjp167, dut_im_yjp167); end else begin $fwrite(tri_report, "Item167 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per167, gol_im_yjp167, dut_im_yjp167); end end

if(col_index>=168) begin if(err_re_per168 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item168 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per168, gol_re_yjp168, dut_re_yjp168); end else begin $fwrite(tri_report, "Item168 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per168, gol_re_yjp168, dut_re_yjp168); end end
if(col_index>=168) begin if(err_im_per168 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item168 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per168, gol_im_yjp168, dut_im_yjp168); end else begin $fwrite(tri_report, "Item168 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per168, gol_im_yjp168, dut_im_yjp168); end end

if(col_index>=169) begin if(err_re_per169 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item169 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per169, gol_re_yjp169, dut_re_yjp169); end else begin $fwrite(tri_report, "Item169 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per169, gol_re_yjp169, dut_re_yjp169); end end
if(col_index>=169) begin if(err_im_per169 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item169 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per169, gol_im_yjp169, dut_im_yjp169); end else begin $fwrite(tri_report, "Item169 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per169, gol_im_yjp169, dut_im_yjp169); end end

if(col_index>=170) begin if(err_re_per170 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item170 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per170, gol_re_yjp170, dut_re_yjp170); end else begin $fwrite(tri_report, "Item170 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per170, gol_re_yjp170, dut_re_yjp170); end end
if(col_index>=170) begin if(err_im_per170 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item170 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per170, gol_im_yjp170, dut_im_yjp170); end else begin $fwrite(tri_report, "Item170 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per170, gol_im_yjp170, dut_im_yjp170); end end

if(col_index>=171) begin if(err_re_per171 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item171 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per171, gol_re_yjp171, dut_re_yjp171); end else begin $fwrite(tri_report, "Item171 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per171, gol_re_yjp171, dut_re_yjp171); end end
if(col_index>=171) begin if(err_im_per171 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item171 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per171, gol_im_yjp171, dut_im_yjp171); end else begin $fwrite(tri_report, "Item171 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per171, gol_im_yjp171, dut_im_yjp171); end end

if(col_index>=172) begin if(err_re_per172 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item172 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per172, gol_re_yjp172, dut_re_yjp172); end else begin $fwrite(tri_report, "Item172 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per172, gol_re_yjp172, dut_re_yjp172); end end
if(col_index>=172) begin if(err_im_per172 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item172 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per172, gol_im_yjp172, dut_im_yjp172); end else begin $fwrite(tri_report, "Item172 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per172, gol_im_yjp172, dut_im_yjp172); end end

if(col_index>=173) begin if(err_re_per173 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item173 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per173, gol_re_yjp173, dut_re_yjp173); end else begin $fwrite(tri_report, "Item173 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per173, gol_re_yjp173, dut_re_yjp173); end end
if(col_index>=173) begin if(err_im_per173 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item173 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per173, gol_im_yjp173, dut_im_yjp173); end else begin $fwrite(tri_report, "Item173 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per173, gol_im_yjp173, dut_im_yjp173); end end

if(col_index>=174) begin if(err_re_per174 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item174 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per174, gol_re_yjp174, dut_re_yjp174); end else begin $fwrite(tri_report, "Item174 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per174, gol_re_yjp174, dut_re_yjp174); end end
if(col_index>=174) begin if(err_im_per174 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item174 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per174, gol_im_yjp174, dut_im_yjp174); end else begin $fwrite(tri_report, "Item174 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per174, gol_im_yjp174, dut_im_yjp174); end end

if(col_index>=175) begin if(err_re_per175 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item175 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per175, gol_re_yjp175, dut_re_yjp175); end else begin $fwrite(tri_report, "Item175 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per175, gol_re_yjp175, dut_re_yjp175); end end
if(col_index>=175) begin if(err_im_per175 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item175 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per175, gol_im_yjp175, dut_im_yjp175); end else begin $fwrite(tri_report, "Item175 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per175, gol_im_yjp175, dut_im_yjp175); end end

if(col_index>=176) begin if(err_re_per176 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item176 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per176, gol_re_yjp176, dut_re_yjp176); end else begin $fwrite(tri_report, "Item176 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per176, gol_re_yjp176, dut_re_yjp176); end end
if(col_index>=176) begin if(err_im_per176 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item176 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per176, gol_im_yjp176, dut_im_yjp176); end else begin $fwrite(tri_report, "Item176 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per176, gol_im_yjp176, dut_im_yjp176); end end

if(col_index>=177) begin if(err_re_per177 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item177 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per177, gol_re_yjp177, dut_re_yjp177); end else begin $fwrite(tri_report, "Item177 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per177, gol_re_yjp177, dut_re_yjp177); end end
if(col_index>=177) begin if(err_im_per177 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item177 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per177, gol_im_yjp177, dut_im_yjp177); end else begin $fwrite(tri_report, "Item177 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per177, gol_im_yjp177, dut_im_yjp177); end end

if(col_index>=178) begin if(err_re_per178 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item178 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per178, gol_re_yjp178, dut_re_yjp178); end else begin $fwrite(tri_report, "Item178 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per178, gol_re_yjp178, dut_re_yjp178); end end
if(col_index>=178) begin if(err_im_per178 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item178 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per178, gol_im_yjp178, dut_im_yjp178); end else begin $fwrite(tri_report, "Item178 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per178, gol_im_yjp178, dut_im_yjp178); end end

if(col_index>=179) begin if(err_re_per179 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item179 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per179, gol_re_yjp179, dut_re_yjp179); end else begin $fwrite(tri_report, "Item179 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per179, gol_re_yjp179, dut_re_yjp179); end end
if(col_index>=179) begin if(err_im_per179 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item179 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per179, gol_im_yjp179, dut_im_yjp179); end else begin $fwrite(tri_report, "Item179 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per179, gol_im_yjp179, dut_im_yjp179); end end

if(col_index>=180) begin if(err_re_per180 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item180 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per180, gol_re_yjp180, dut_re_yjp180); end else begin $fwrite(tri_report, "Item180 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per180, gol_re_yjp180, dut_re_yjp180); end end
if(col_index>=180) begin if(err_im_per180 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item180 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per180, gol_im_yjp180, dut_im_yjp180); end else begin $fwrite(tri_report, "Item180 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per180, gol_im_yjp180, dut_im_yjp180); end end

if(col_index>=181) begin if(err_re_per181 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item181 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per181, gol_re_yjp181, dut_re_yjp181); end else begin $fwrite(tri_report, "Item181 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per181, gol_re_yjp181, dut_re_yjp181); end end
if(col_index>=181) begin if(err_im_per181 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item181 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per181, gol_im_yjp181, dut_im_yjp181); end else begin $fwrite(tri_report, "Item181 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per181, gol_im_yjp181, dut_im_yjp181); end end

if(col_index>=182) begin if(err_re_per182 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item182 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per182, gol_re_yjp182, dut_re_yjp182); end else begin $fwrite(tri_report, "Item182 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per182, gol_re_yjp182, dut_re_yjp182); end end
if(col_index>=182) begin if(err_im_per182 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item182 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per182, gol_im_yjp182, dut_im_yjp182); end else begin $fwrite(tri_report, "Item182 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per182, gol_im_yjp182, dut_im_yjp182); end end

if(col_index>=183) begin if(err_re_per183 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item183 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per183, gol_re_yjp183, dut_re_yjp183); end else begin $fwrite(tri_report, "Item183 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per183, gol_re_yjp183, dut_re_yjp183); end end
if(col_index>=183) begin if(err_im_per183 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item183 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per183, gol_im_yjp183, dut_im_yjp183); end else begin $fwrite(tri_report, "Item183 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per183, gol_im_yjp183, dut_im_yjp183); end end

if(col_index>=184) begin if(err_re_per184 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item184 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per184, gol_re_yjp184, dut_re_yjp184); end else begin $fwrite(tri_report, "Item184 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per184, gol_re_yjp184, dut_re_yjp184); end end
if(col_index>=184) begin if(err_im_per184 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item184 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per184, gol_im_yjp184, dut_im_yjp184); end else begin $fwrite(tri_report, "Item184 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per184, gol_im_yjp184, dut_im_yjp184); end end

if(col_index>=185) begin if(err_re_per185 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item185 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per185, gol_re_yjp185, dut_re_yjp185); end else begin $fwrite(tri_report, "Item185 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per185, gol_re_yjp185, dut_re_yjp185); end end
if(col_index>=185) begin if(err_im_per185 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item185 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per185, gol_im_yjp185, dut_im_yjp185); end else begin $fwrite(tri_report, "Item185 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per185, gol_im_yjp185, dut_im_yjp185); end end

if(col_index>=186) begin if(err_re_per186 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item186 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per186, gol_re_yjp186, dut_re_yjp186); end else begin $fwrite(tri_report, "Item186 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per186, gol_re_yjp186, dut_re_yjp186); end end
if(col_index>=186) begin if(err_im_per186 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item186 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per186, gol_im_yjp186, dut_im_yjp186); end else begin $fwrite(tri_report, "Item186 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per186, gol_im_yjp186, dut_im_yjp186); end end

if(col_index>=187) begin if(err_re_per187 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item187 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per187, gol_re_yjp187, dut_re_yjp187); end else begin $fwrite(tri_report, "Item187 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per187, gol_re_yjp187, dut_re_yjp187); end end
if(col_index>=187) begin if(err_im_per187 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item187 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per187, gol_im_yjp187, dut_im_yjp187); end else begin $fwrite(tri_report, "Item187 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per187, gol_im_yjp187, dut_im_yjp187); end end

if(col_index>=188) begin if(err_re_per188 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item188 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per188, gol_re_yjp188, dut_re_yjp188); end else begin $fwrite(tri_report, "Item188 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per188, gol_re_yjp188, dut_re_yjp188); end end
if(col_index>=188) begin if(err_im_per188 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item188 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per188, gol_im_yjp188, dut_im_yjp188); end else begin $fwrite(tri_report, "Item188 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per188, gol_im_yjp188, dut_im_yjp188); end end

if(col_index>=189) begin if(err_re_per189 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item189 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per189, gol_re_yjp189, dut_re_yjp189); end else begin $fwrite(tri_report, "Item189 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per189, gol_re_yjp189, dut_re_yjp189); end end
if(col_index>=189) begin if(err_im_per189 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item189 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per189, gol_im_yjp189, dut_im_yjp189); end else begin $fwrite(tri_report, "Item189 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per189, gol_im_yjp189, dut_im_yjp189); end end

if(col_index>=190) begin if(err_re_per190 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item190 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per190, gol_re_yjp190, dut_re_yjp190); end else begin $fwrite(tri_report, "Item190 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per190, gol_re_yjp190, dut_re_yjp190); end end
if(col_index>=190) begin if(err_im_per190 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item190 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per190, gol_im_yjp190, dut_im_yjp190); end else begin $fwrite(tri_report, "Item190 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per190, gol_im_yjp190, dut_im_yjp190); end end

if(col_index>=191) begin if(err_re_per191 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item191 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per191, gol_re_yjp191, dut_re_yjp191); end else begin $fwrite(tri_report, "Item191 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per191, gol_re_yjp191, dut_re_yjp191); end end
if(col_index>=191) begin if(err_im_per191 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item191 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per191, gol_im_yjp191, dut_im_yjp191); end else begin $fwrite(tri_report, "Item191 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per191, gol_im_yjp191, dut_im_yjp191); end end

if(col_index>=192) begin if(err_re_per192 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item192 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per192, gol_re_yjp192, dut_re_yjp192); end else begin $fwrite(tri_report, "Item192 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per192, gol_re_yjp192, dut_re_yjp192); end end
if(col_index>=192) begin if(err_im_per192 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item192 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per192, gol_im_yjp192, dut_im_yjp192); end else begin $fwrite(tri_report, "Item192 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per192, gol_im_yjp192, dut_im_yjp192); end end

if(col_index>=193) begin if(err_re_per193 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item193 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per193, gol_re_yjp193, dut_re_yjp193); end else begin $fwrite(tri_report, "Item193 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per193, gol_re_yjp193, dut_re_yjp193); end end
if(col_index>=193) begin if(err_im_per193 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item193 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per193, gol_im_yjp193, dut_im_yjp193); end else begin $fwrite(tri_report, "Item193 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per193, gol_im_yjp193, dut_im_yjp193); end end

if(col_index>=194) begin if(err_re_per194 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item194 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per194, gol_re_yjp194, dut_re_yjp194); end else begin $fwrite(tri_report, "Item194 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per194, gol_re_yjp194, dut_re_yjp194); end end
if(col_index>=194) begin if(err_im_per194 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item194 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per194, gol_im_yjp194, dut_im_yjp194); end else begin $fwrite(tri_report, "Item194 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per194, gol_im_yjp194, dut_im_yjp194); end end

if(col_index>=195) begin if(err_re_per195 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item195 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per195, gol_re_yjp195, dut_re_yjp195); end else begin $fwrite(tri_report, "Item195 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per195, gol_re_yjp195, dut_re_yjp195); end end
if(col_index>=195) begin if(err_im_per195 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item195 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per195, gol_im_yjp195, dut_im_yjp195); end else begin $fwrite(tri_report, "Item195 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per195, gol_im_yjp195, dut_im_yjp195); end end

if(col_index>=196) begin if(err_re_per196 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item196 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per196, gol_re_yjp196, dut_re_yjp196); end else begin $fwrite(tri_report, "Item196 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per196, gol_re_yjp196, dut_re_yjp196); end end
if(col_index>=196) begin if(err_im_per196 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item196 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per196, gol_im_yjp196, dut_im_yjp196); end else begin $fwrite(tri_report, "Item196 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per196, gol_im_yjp196, dut_im_yjp196); end end

if(col_index>=197) begin if(err_re_per197 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item197 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per197, gol_re_yjp197, dut_re_yjp197); end else begin $fwrite(tri_report, "Item197 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per197, gol_re_yjp197, dut_re_yjp197); end end
if(col_index>=197) begin if(err_im_per197 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item197 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per197, gol_im_yjp197, dut_im_yjp197); end else begin $fwrite(tri_report, "Item197 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per197, gol_im_yjp197, dut_im_yjp197); end end

if(col_index>=198) begin if(err_re_per198 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item198 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per198, gol_re_yjp198, dut_re_yjp198); end else begin $fwrite(tri_report, "Item198 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per198, gol_re_yjp198, dut_re_yjp198); end end
if(col_index>=198) begin if(err_im_per198 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item198 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per198, gol_im_yjp198, dut_im_yjp198); end else begin $fwrite(tri_report, "Item198 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per198, gol_im_yjp198, dut_im_yjp198); end end

if(col_index>=199) begin if(err_re_per199 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item199 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per199, gol_re_yjp199, dut_re_yjp199); end else begin $fwrite(tri_report, "Item199 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per199, gol_re_yjp199, dut_re_yjp199); end end
if(col_index>=199) begin if(err_im_per199 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item199 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per199, gol_im_yjp199, dut_im_yjp199); end else begin $fwrite(tri_report, "Item199 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per199, gol_im_yjp199, dut_im_yjp199); end end

if(col_index>=200) begin if(err_re_per200 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item200 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per200, gol_re_yjp200, dut_re_yjp200); end else begin $fwrite(tri_report, "Item200 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per200, gol_re_yjp200, dut_re_yjp200); end end
if(col_index>=200) begin if(err_im_per200 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item200 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per200, gol_im_yjp200, dut_im_yjp200); end else begin $fwrite(tri_report, "Item200 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per200, gol_im_yjp200, dut_im_yjp200); end end

if(col_index>=201) begin if(err_re_per201 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item201 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per201, gol_re_yjp201, dut_re_yjp201); end else begin $fwrite(tri_report, "Item201 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per201, gol_re_yjp201, dut_re_yjp201); end end
if(col_index>=201) begin if(err_im_per201 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item201 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per201, gol_im_yjp201, dut_im_yjp201); end else begin $fwrite(tri_report, "Item201 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per201, gol_im_yjp201, dut_im_yjp201); end end

if(col_index>=202) begin if(err_re_per202 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item202 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per202, gol_re_yjp202, dut_re_yjp202); end else begin $fwrite(tri_report, "Item202 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per202, gol_re_yjp202, dut_re_yjp202); end end
if(col_index>=202) begin if(err_im_per202 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item202 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per202, gol_im_yjp202, dut_im_yjp202); end else begin $fwrite(tri_report, "Item202 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per202, gol_im_yjp202, dut_im_yjp202); end end

if(col_index>=203) begin if(err_re_per203 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item203 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per203, gol_re_yjp203, dut_re_yjp203); end else begin $fwrite(tri_report, "Item203 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per203, gol_re_yjp203, dut_re_yjp203); end end
if(col_index>=203) begin if(err_im_per203 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item203 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per203, gol_im_yjp203, dut_im_yjp203); end else begin $fwrite(tri_report, "Item203 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per203, gol_im_yjp203, dut_im_yjp203); end end

if(col_index>=204) begin if(err_re_per204 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item204 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per204, gol_re_yjp204, dut_re_yjp204); end else begin $fwrite(tri_report, "Item204 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per204, gol_re_yjp204, dut_re_yjp204); end end
if(col_index>=204) begin if(err_im_per204 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item204 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per204, gol_im_yjp204, dut_im_yjp204); end else begin $fwrite(tri_report, "Item204 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per204, gol_im_yjp204, dut_im_yjp204); end end

if(col_index>=205) begin if(err_re_per205 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item205 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per205, gol_re_yjp205, dut_re_yjp205); end else begin $fwrite(tri_report, "Item205 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per205, gol_re_yjp205, dut_re_yjp205); end end
if(col_index>=205) begin if(err_im_per205 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item205 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per205, gol_im_yjp205, dut_im_yjp205); end else begin $fwrite(tri_report, "Item205 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per205, gol_im_yjp205, dut_im_yjp205); end end

if(col_index>=206) begin if(err_re_per206 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item206 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per206, gol_re_yjp206, dut_re_yjp206); end else begin $fwrite(tri_report, "Item206 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per206, gol_re_yjp206, dut_re_yjp206); end end
if(col_index>=206) begin if(err_im_per206 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item206 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per206, gol_im_yjp206, dut_im_yjp206); end else begin $fwrite(tri_report, "Item206 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per206, gol_im_yjp206, dut_im_yjp206); end end

if(col_index>=207) begin if(err_re_per207 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item207 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per207, gol_re_yjp207, dut_re_yjp207); end else begin $fwrite(tri_report, "Item207 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per207, gol_re_yjp207, dut_re_yjp207); end end
if(col_index>=207) begin if(err_im_per207 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item207 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per207, gol_im_yjp207, dut_im_yjp207); end else begin $fwrite(tri_report, "Item207 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per207, gol_im_yjp207, dut_im_yjp207); end end

if(col_index>=208) begin if(err_re_per208 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item208 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per208, gol_re_yjp208, dut_re_yjp208); end else begin $fwrite(tri_report, "Item208 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per208, gol_re_yjp208, dut_re_yjp208); end end
if(col_index>=208) begin if(err_im_per208 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item208 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per208, gol_im_yjp208, dut_im_yjp208); end else begin $fwrite(tri_report, "Item208 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per208, gol_im_yjp208, dut_im_yjp208); end end

if(col_index>=209) begin if(err_re_per209 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item209 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per209, gol_re_yjp209, dut_re_yjp209); end else begin $fwrite(tri_report, "Item209 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per209, gol_re_yjp209, dut_re_yjp209); end end
if(col_index>=209) begin if(err_im_per209 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item209 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per209, gol_im_yjp209, dut_im_yjp209); end else begin $fwrite(tri_report, "Item209 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per209, gol_im_yjp209, dut_im_yjp209); end end

if(col_index>=210) begin if(err_re_per210 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item210 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per210, gol_re_yjp210, dut_re_yjp210); end else begin $fwrite(tri_report, "Item210 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per210, gol_re_yjp210, dut_re_yjp210); end end
if(col_index>=210) begin if(err_im_per210 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item210 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per210, gol_im_yjp210, dut_im_yjp210); end else begin $fwrite(tri_report, "Item210 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per210, gol_im_yjp210, dut_im_yjp210); end end

if(col_index>=211) begin if(err_re_per211 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item211 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per211, gol_re_yjp211, dut_re_yjp211); end else begin $fwrite(tri_report, "Item211 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per211, gol_re_yjp211, dut_re_yjp211); end end
if(col_index>=211) begin if(err_im_per211 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item211 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per211, gol_im_yjp211, dut_im_yjp211); end else begin $fwrite(tri_report, "Item211 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per211, gol_im_yjp211, dut_im_yjp211); end end

if(col_index>=212) begin if(err_re_per212 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item212 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per212, gol_re_yjp212, dut_re_yjp212); end else begin $fwrite(tri_report, "Item212 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per212, gol_re_yjp212, dut_re_yjp212); end end
if(col_index>=212) begin if(err_im_per212 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item212 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per212, gol_im_yjp212, dut_im_yjp212); end else begin $fwrite(tri_report, "Item212 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per212, gol_im_yjp212, dut_im_yjp212); end end

if(col_index>=213) begin if(err_re_per213 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item213 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per213, gol_re_yjp213, dut_re_yjp213); end else begin $fwrite(tri_report, "Item213 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per213, gol_re_yjp213, dut_re_yjp213); end end
if(col_index>=213) begin if(err_im_per213 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item213 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per213, gol_im_yjp213, dut_im_yjp213); end else begin $fwrite(tri_report, "Item213 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per213, gol_im_yjp213, dut_im_yjp213); end end

if(col_index>=214) begin if(err_re_per214 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item214 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per214, gol_re_yjp214, dut_re_yjp214); end else begin $fwrite(tri_report, "Item214 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per214, gol_re_yjp214, dut_re_yjp214); end end
if(col_index>=214) begin if(err_im_per214 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item214 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per214, gol_im_yjp214, dut_im_yjp214); end else begin $fwrite(tri_report, "Item214 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per214, gol_im_yjp214, dut_im_yjp214); end end

if(col_index>=215) begin if(err_re_per215 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item215 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per215, gol_re_yjp215, dut_re_yjp215); end else begin $fwrite(tri_report, "Item215 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per215, gol_re_yjp215, dut_re_yjp215); end end
if(col_index>=215) begin if(err_im_per215 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item215 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per215, gol_im_yjp215, dut_im_yjp215); end else begin $fwrite(tri_report, "Item215 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per215, gol_im_yjp215, dut_im_yjp215); end end

if(col_index>=216) begin if(err_re_per216 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item216 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per216, gol_re_yjp216, dut_re_yjp216); end else begin $fwrite(tri_report, "Item216 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per216, gol_re_yjp216, dut_re_yjp216); end end
if(col_index>=216) begin if(err_im_per216 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item216 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per216, gol_im_yjp216, dut_im_yjp216); end else begin $fwrite(tri_report, "Item216 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per216, gol_im_yjp216, dut_im_yjp216); end end

if(col_index>=217) begin if(err_re_per217 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item217 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per217, gol_re_yjp217, dut_re_yjp217); end else begin $fwrite(tri_report, "Item217 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per217, gol_re_yjp217, dut_re_yjp217); end end
if(col_index>=217) begin if(err_im_per217 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item217 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per217, gol_im_yjp217, dut_im_yjp217); end else begin $fwrite(tri_report, "Item217 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per217, gol_im_yjp217, dut_im_yjp217); end end

if(col_index>=218) begin if(err_re_per218 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item218 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per218, gol_re_yjp218, dut_re_yjp218); end else begin $fwrite(tri_report, "Item218 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per218, gol_re_yjp218, dut_re_yjp218); end end
if(col_index>=218) begin if(err_im_per218 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item218 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per218, gol_im_yjp218, dut_im_yjp218); end else begin $fwrite(tri_report, "Item218 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per218, gol_im_yjp218, dut_im_yjp218); end end

if(col_index>=219) begin if(err_re_per219 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item219 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per219, gol_re_yjp219, dut_re_yjp219); end else begin $fwrite(tri_report, "Item219 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per219, gol_re_yjp219, dut_re_yjp219); end end
if(col_index>=219) begin if(err_im_per219 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item219 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per219, gol_im_yjp219, dut_im_yjp219); end else begin $fwrite(tri_report, "Item219 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per219, gol_im_yjp219, dut_im_yjp219); end end

if(col_index>=220) begin if(err_re_per220 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item220 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per220, gol_re_yjp220, dut_re_yjp220); end else begin $fwrite(tri_report, "Item220 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per220, gol_re_yjp220, dut_re_yjp220); end end
if(col_index>=220) begin if(err_im_per220 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item220 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per220, gol_im_yjp220, dut_im_yjp220); end else begin $fwrite(tri_report, "Item220 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per220, gol_im_yjp220, dut_im_yjp220); end end

if(col_index>=221) begin if(err_re_per221 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item221 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per221, gol_re_yjp221, dut_re_yjp221); end else begin $fwrite(tri_report, "Item221 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per221, gol_re_yjp221, dut_re_yjp221); end end
if(col_index>=221) begin if(err_im_per221 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item221 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per221, gol_im_yjp221, dut_im_yjp221); end else begin $fwrite(tri_report, "Item221 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per221, gol_im_yjp221, dut_im_yjp221); end end

if(col_index>=222) begin if(err_re_per222 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item222 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per222, gol_re_yjp222, dut_re_yjp222); end else begin $fwrite(tri_report, "Item222 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per222, gol_re_yjp222, dut_re_yjp222); end end
if(col_index>=222) begin if(err_im_per222 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item222 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per222, gol_im_yjp222, dut_im_yjp222); end else begin $fwrite(tri_report, "Item222 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per222, gol_im_yjp222, dut_im_yjp222); end end

if(col_index>=223) begin if(err_re_per223 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item223 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per223, gol_re_yjp223, dut_re_yjp223); end else begin $fwrite(tri_report, "Item223 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per223, gol_re_yjp223, dut_re_yjp223); end end
if(col_index>=223) begin if(err_im_per223 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item223 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per223, gol_im_yjp223, dut_im_yjp223); end else begin $fwrite(tri_report, "Item223 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per223, gol_im_yjp223, dut_im_yjp223); end end

if(col_index>=224) begin if(err_re_per224 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item224 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per224, gol_re_yjp224, dut_re_yjp224); end else begin $fwrite(tri_report, "Item224 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per224, gol_re_yjp224, dut_re_yjp224); end end
if(col_index>=224) begin if(err_im_per224 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item224 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per224, gol_im_yjp224, dut_im_yjp224); end else begin $fwrite(tri_report, "Item224 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per224, gol_im_yjp224, dut_im_yjp224); end end

if(col_index>=225) begin if(err_re_per225 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item225 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per225, gol_re_yjp225, dut_re_yjp225); end else begin $fwrite(tri_report, "Item225 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per225, gol_re_yjp225, dut_re_yjp225); end end
if(col_index>=225) begin if(err_im_per225 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item225 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per225, gol_im_yjp225, dut_im_yjp225); end else begin $fwrite(tri_report, "Item225 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per225, gol_im_yjp225, dut_im_yjp225); end end

if(col_index>=226) begin if(err_re_per226 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item226 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per226, gol_re_yjp226, dut_re_yjp226); end else begin $fwrite(tri_report, "Item226 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per226, gol_re_yjp226, dut_re_yjp226); end end
if(col_index>=226) begin if(err_im_per226 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item226 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per226, gol_im_yjp226, dut_im_yjp226); end else begin $fwrite(tri_report, "Item226 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per226, gol_im_yjp226, dut_im_yjp226); end end

if(col_index>=227) begin if(err_re_per227 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item227 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per227, gol_re_yjp227, dut_re_yjp227); end else begin $fwrite(tri_report, "Item227 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per227, gol_re_yjp227, dut_re_yjp227); end end
if(col_index>=227) begin if(err_im_per227 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item227 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per227, gol_im_yjp227, dut_im_yjp227); end else begin $fwrite(tri_report, "Item227 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per227, gol_im_yjp227, dut_im_yjp227); end end

if(col_index>=228) begin if(err_re_per228 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item228 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per228, gol_re_yjp228, dut_re_yjp228); end else begin $fwrite(tri_report, "Item228 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per228, gol_re_yjp228, dut_re_yjp228); end end
if(col_index>=228) begin if(err_im_per228 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item228 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per228, gol_im_yjp228, dut_im_yjp228); end else begin $fwrite(tri_report, "Item228 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per228, gol_im_yjp228, dut_im_yjp228); end end

if(col_index>=229) begin if(err_re_per229 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item229 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per229, gol_re_yjp229, dut_re_yjp229); end else begin $fwrite(tri_report, "Item229 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per229, gol_re_yjp229, dut_re_yjp229); end end
if(col_index>=229) begin if(err_im_per229 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item229 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per229, gol_im_yjp229, dut_im_yjp229); end else begin $fwrite(tri_report, "Item229 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per229, gol_im_yjp229, dut_im_yjp229); end end

if(col_index>=230) begin if(err_re_per230 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item230 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per230, gol_re_yjp230, dut_re_yjp230); end else begin $fwrite(tri_report, "Item230 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per230, gol_re_yjp230, dut_re_yjp230); end end
if(col_index>=230) begin if(err_im_per230 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item230 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per230, gol_im_yjp230, dut_im_yjp230); end else begin $fwrite(tri_report, "Item230 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per230, gol_im_yjp230, dut_im_yjp230); end end

if(col_index>=231) begin if(err_re_per231 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item231 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per231, gol_re_yjp231, dut_re_yjp231); end else begin $fwrite(tri_report, "Item231 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per231, gol_re_yjp231, dut_re_yjp231); end end
if(col_index>=231) begin if(err_im_per231 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item231 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per231, gol_im_yjp231, dut_im_yjp231); end else begin $fwrite(tri_report, "Item231 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per231, gol_im_yjp231, dut_im_yjp231); end end

if(col_index>=232) begin if(err_re_per232 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item232 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per232, gol_re_yjp232, dut_re_yjp232); end else begin $fwrite(tri_report, "Item232 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per232, gol_re_yjp232, dut_re_yjp232); end end
if(col_index>=232) begin if(err_im_per232 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item232 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per232, gol_im_yjp232, dut_im_yjp232); end else begin $fwrite(tri_report, "Item232 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per232, gol_im_yjp232, dut_im_yjp232); end end

if(col_index>=233) begin if(err_re_per233 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item233 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per233, gol_re_yjp233, dut_re_yjp233); end else begin $fwrite(tri_report, "Item233 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per233, gol_re_yjp233, dut_re_yjp233); end end
if(col_index>=233) begin if(err_im_per233 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item233 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per233, gol_im_yjp233, dut_im_yjp233); end else begin $fwrite(tri_report, "Item233 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per233, gol_im_yjp233, dut_im_yjp233); end end

if(col_index>=234) begin if(err_re_per234 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item234 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per234, gol_re_yjp234, dut_re_yjp234); end else begin $fwrite(tri_report, "Item234 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per234, gol_re_yjp234, dut_re_yjp234); end end
if(col_index>=234) begin if(err_im_per234 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item234 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per234, gol_im_yjp234, dut_im_yjp234); end else begin $fwrite(tri_report, "Item234 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per234, gol_im_yjp234, dut_im_yjp234); end end

if(col_index>=235) begin if(err_re_per235 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item235 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per235, gol_re_yjp235, dut_re_yjp235); end else begin $fwrite(tri_report, "Item235 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per235, gol_re_yjp235, dut_re_yjp235); end end
if(col_index>=235) begin if(err_im_per235 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item235 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per235, gol_im_yjp235, dut_im_yjp235); end else begin $fwrite(tri_report, "Item235 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per235, gol_im_yjp235, dut_im_yjp235); end end

if(col_index>=236) begin if(err_re_per236 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item236 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per236, gol_re_yjp236, dut_re_yjp236); end else begin $fwrite(tri_report, "Item236 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per236, gol_re_yjp236, dut_re_yjp236); end end
if(col_index>=236) begin if(err_im_per236 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item236 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per236, gol_im_yjp236, dut_im_yjp236); end else begin $fwrite(tri_report, "Item236 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per236, gol_im_yjp236, dut_im_yjp236); end end

if(col_index>=237) begin if(err_re_per237 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item237 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per237, gol_re_yjp237, dut_re_yjp237); end else begin $fwrite(tri_report, "Item237 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per237, gol_re_yjp237, dut_re_yjp237); end end
if(col_index>=237) begin if(err_im_per237 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item237 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per237, gol_im_yjp237, dut_im_yjp237); end else begin $fwrite(tri_report, "Item237 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per237, gol_im_yjp237, dut_im_yjp237); end end

if(col_index>=238) begin if(err_re_per238 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item238 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per238, gol_re_yjp238, dut_re_yjp238); end else begin $fwrite(tri_report, "Item238 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per238, gol_re_yjp238, dut_re_yjp238); end end
if(col_index>=238) begin if(err_im_per238 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item238 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per238, gol_im_yjp238, dut_im_yjp238); end else begin $fwrite(tri_report, "Item238 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per238, gol_im_yjp238, dut_im_yjp238); end end

if(col_index>=239) begin if(err_re_per239 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item239 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per239, gol_re_yjp239, dut_re_yjp239); end else begin $fwrite(tri_report, "Item239 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per239, gol_re_yjp239, dut_re_yjp239); end end
if(col_index>=239) begin if(err_im_per239 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item239 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per239, gol_im_yjp239, dut_im_yjp239); end else begin $fwrite(tri_report, "Item239 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per239, gol_im_yjp239, dut_im_yjp239); end end

if(col_index>=240) begin if(err_re_per240 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item240 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per240, gol_re_yjp240, dut_re_yjp240); end else begin $fwrite(tri_report, "Item240 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per240, gol_re_yjp240, dut_re_yjp240); end end
if(col_index>=240) begin if(err_im_per240 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item240 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per240, gol_im_yjp240, dut_im_yjp240); end else begin $fwrite(tri_report, "Item240 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per240, gol_im_yjp240, dut_im_yjp240); end end

if(col_index>=241) begin if(err_re_per241 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item241 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per241, gol_re_yjp241, dut_re_yjp241); end else begin $fwrite(tri_report, "Item241 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per241, gol_re_yjp241, dut_re_yjp241); end end
if(col_index>=241) begin if(err_im_per241 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item241 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per241, gol_im_yjp241, dut_im_yjp241); end else begin $fwrite(tri_report, "Item241 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per241, gol_im_yjp241, dut_im_yjp241); end end

if(col_index>=242) begin if(err_re_per242 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item242 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per242, gol_re_yjp242, dut_re_yjp242); end else begin $fwrite(tri_report, "Item242 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per242, gol_re_yjp242, dut_re_yjp242); end end
if(col_index>=242) begin if(err_im_per242 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item242 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per242, gol_im_yjp242, dut_im_yjp242); end else begin $fwrite(tri_report, "Item242 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per242, gol_im_yjp242, dut_im_yjp242); end end

if(col_index>=243) begin if(err_re_per243 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item243 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per243, gol_re_yjp243, dut_re_yjp243); end else begin $fwrite(tri_report, "Item243 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per243, gol_re_yjp243, dut_re_yjp243); end end
if(col_index>=243) begin if(err_im_per243 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item243 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per243, gol_im_yjp243, dut_im_yjp243); end else begin $fwrite(tri_report, "Item243 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per243, gol_im_yjp243, dut_im_yjp243); end end

if(col_index>=244) begin if(err_re_per244 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item244 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per244, gol_re_yjp244, dut_re_yjp244); end else begin $fwrite(tri_report, "Item244 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per244, gol_re_yjp244, dut_re_yjp244); end end
if(col_index>=244) begin if(err_im_per244 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item244 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per244, gol_im_yjp244, dut_im_yjp244); end else begin $fwrite(tri_report, "Item244 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per244, gol_im_yjp244, dut_im_yjp244); end end

if(col_index>=245) begin if(err_re_per245 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item245 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per245, gol_re_yjp245, dut_re_yjp245); end else begin $fwrite(tri_report, "Item245 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per245, gol_re_yjp245, dut_re_yjp245); end end
if(col_index>=245) begin if(err_im_per245 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item245 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per245, gol_im_yjp245, dut_im_yjp245); end else begin $fwrite(tri_report, "Item245 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per245, gol_im_yjp245, dut_im_yjp245); end end

if(col_index>=246) begin if(err_re_per246 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item246 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per246, gol_re_yjp246, dut_re_yjp246); end else begin $fwrite(tri_report, "Item246 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per246, gol_re_yjp246, dut_re_yjp246); end end
if(col_index>=246) begin if(err_im_per246 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item246 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per246, gol_im_yjp246, dut_im_yjp246); end else begin $fwrite(tri_report, "Item246 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per246, gol_im_yjp246, dut_im_yjp246); end end

if(col_index>=247) begin if(err_re_per247 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item247 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per247, gol_re_yjp247, dut_re_yjp247); end else begin $fwrite(tri_report, "Item247 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per247, gol_re_yjp247, dut_re_yjp247); end end
if(col_index>=247) begin if(err_im_per247 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item247 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per247, gol_im_yjp247, dut_im_yjp247); end else begin $fwrite(tri_report, "Item247 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per247, gol_im_yjp247, dut_im_yjp247); end end

if(col_index>=248) begin if(err_re_per248 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item248 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per248, gol_re_yjp248, dut_re_yjp248); end else begin $fwrite(tri_report, "Item248 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per248, gol_re_yjp248, dut_re_yjp248); end end
if(col_index>=248) begin if(err_im_per248 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item248 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per248, gol_im_yjp248, dut_im_yjp248); end else begin $fwrite(tri_report, "Item248 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per248, gol_im_yjp248, dut_im_yjp248); end end

if(col_index>=249) begin if(err_re_per249 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item249 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per249, gol_re_yjp249, dut_re_yjp249); end else begin $fwrite(tri_report, "Item249 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per249, gol_re_yjp249, dut_re_yjp249); end end
if(col_index>=249) begin if(err_im_per249 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item249 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per249, gol_im_yjp249, dut_im_yjp249); end else begin $fwrite(tri_report, "Item249 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per249, gol_im_yjp249, dut_im_yjp249); end end

if(col_index>=250) begin if(err_re_per250 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item250 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per250, gol_re_yjp250, dut_re_yjp250); end else begin $fwrite(tri_report, "Item250 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per250, gol_re_yjp250, dut_re_yjp250); end end
if(col_index>=250) begin if(err_im_per250 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item250 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per250, gol_im_yjp250, dut_im_yjp250); end else begin $fwrite(tri_report, "Item250 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per250, gol_im_yjp250, dut_im_yjp250); end end

if(col_index>=251) begin if(err_re_per251 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item251 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per251, gol_re_yjp251, dut_re_yjp251); end else begin $fwrite(tri_report, "Item251 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per251, gol_re_yjp251, dut_re_yjp251); end end
if(col_index>=251) begin if(err_im_per251 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item251 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per251, gol_im_yjp251, dut_im_yjp251); end else begin $fwrite(tri_report, "Item251 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per251, gol_im_yjp251, dut_im_yjp251); end end

if(col_index>=252) begin if(err_re_per252 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item252 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per252, gol_re_yjp252, dut_re_yjp252); end else begin $fwrite(tri_report, "Item252 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per252, gol_re_yjp252, dut_re_yjp252); end end
if(col_index>=252) begin if(err_im_per252 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item252 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per252, gol_im_yjp252, dut_im_yjp252); end else begin $fwrite(tri_report, "Item252 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per252, gol_im_yjp252, dut_im_yjp252); end end

if(col_index>=253) begin if(err_re_per253 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item253 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per253, gol_re_yjp253, dut_re_yjp253); end else begin $fwrite(tri_report, "Item253 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per253, gol_re_yjp253, dut_re_yjp253); end end
if(col_index>=253) begin if(err_im_per253 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item253 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per253, gol_im_yjp253, dut_im_yjp253); end else begin $fwrite(tri_report, "Item253 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per253, gol_im_yjp253, dut_im_yjp253); end end

if(col_index>=254) begin if(err_re_per254 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item254 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per254, gol_re_yjp254, dut_re_yjp254); end else begin $fwrite(tri_report, "Item254 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per254, gol_re_yjp254, dut_re_yjp254); end end
if(col_index>=254) begin if(err_im_per254 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item254 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per254, gol_im_yjp254, dut_im_yjp254); end else begin $fwrite(tri_report, "Item254 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per254, gol_im_yjp254, dut_im_yjp254); end end

if(col_index>=255) begin if(err_re_per255 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item255 Re Comp Pass! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per255, gol_re_yjp255, dut_re_yjp255); end else begin $fwrite(tri_report, "Item255 Re  Comp FAIL! error real percent: %f%%, golden real result: %f, dut real result: %f\n", err_re_per255, gol_re_yjp255, dut_re_yjp255); end end
if(col_index>=255) begin if(err_im_per255 <= `ERROR_THRESHOLD) begin $fwrite(tri_report, "Item255 Im  Comp Pass! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per255, gol_im_yjp255, dut_im_yjp255); end else begin $fwrite(tri_report, "Item255 Im Comp FAIL! error imaginary percent: %f%%, golden imaginary result: %f, dut imaginary result: %f\n", err_im_per255, gol_im_yjp255, dut_im_yjp255); end end

`endif

